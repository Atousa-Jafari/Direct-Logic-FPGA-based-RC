`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 03/04/2024 09:10:17 AM
// Design Name:
// Module Name: EchoStateNetwork
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

(* use_dsp="yes" *)module ESN_Generator_V2(
    input clk,
    input signed [7:0] input_data,
    output wire signed [31:0] output_data
);
parameter num_reservoir_neurons = 200;

// Input layer
reg signed [7:0] input_weight [0: num_reservoir_neurons-1];
initial {
input_weight[0],
input_weight[1],
input_weight[2],
input_weight[3],
input_weight[4],
input_weight[5],
input_weight[6],
input_weight[7],
input_weight[8],
input_weight[9],
input_weight[10],
input_weight[11],
input_weight[12],
input_weight[13],
input_weight[14],
input_weight[15],
input_weight[16],
input_weight[17],
input_weight[18],
input_weight[19],
input_weight[20],
input_weight[21],
input_weight[22],
input_weight[23],
input_weight[24],
input_weight[25],
input_weight[26],
input_weight[27],
input_weight[28],
input_weight[29],
input_weight[30],
input_weight[31],
input_weight[32],
input_weight[33],
input_weight[34],
input_weight[35],
input_weight[36],
input_weight[37],
input_weight[38],
input_weight[39],
input_weight[40],
input_weight[41],
input_weight[42],
input_weight[43],
input_weight[44],
input_weight[45],
input_weight[46],
input_weight[47],
input_weight[48],
input_weight[49],
input_weight[50],
input_weight[51],
input_weight[52],
input_weight[53],
input_weight[54],
input_weight[55],
input_weight[56],
input_weight[57],
input_weight[58],
input_weight[59],
input_weight[60],
input_weight[61],
input_weight[62],
input_weight[63],
input_weight[64],
input_weight[65],
input_weight[66],
input_weight[67],
input_weight[68],
input_weight[69],
input_weight[70],
input_weight[71],
input_weight[72],
input_weight[73],
input_weight[74],
input_weight[75],
input_weight[76],
input_weight[77],
input_weight[78],
input_weight[79],
input_weight[80],
input_weight[81],
input_weight[82],
input_weight[83],
input_weight[84],
input_weight[85],
input_weight[86],
input_weight[87],
input_weight[88],
input_weight[89],
input_weight[90],
input_weight[91],
input_weight[92],
input_weight[93],
input_weight[94],
input_weight[95],
input_weight[96],
input_weight[97],
input_weight[98],
input_weight[99],
input_weight[100],
input_weight[101],
input_weight[102],
input_weight[103],
input_weight[104],
input_weight[105],
input_weight[106],
input_weight[107],
input_weight[108],
input_weight[109],
input_weight[110],
input_weight[111],
input_weight[112],
input_weight[113],
input_weight[114],
input_weight[115],
input_weight[116],
input_weight[117],
input_weight[118],
input_weight[119],
input_weight[120],
input_weight[121],
input_weight[122],
input_weight[123],
input_weight[124],
input_weight[125],
input_weight[126],
input_weight[127],
input_weight[128],
input_weight[129],
input_weight[130],
input_weight[131],
input_weight[132],
input_weight[133],
input_weight[134],
input_weight[135],
input_weight[136],
input_weight[137],
input_weight[138],
input_weight[139],
input_weight[140],
input_weight[141],
input_weight[142],
input_weight[143],
input_weight[144],
input_weight[145],
input_weight[146],
input_weight[147],
input_weight[148],
input_weight[149],
input_weight[150],
input_weight[151],
input_weight[152],
input_weight[153],
input_weight[154],
input_weight[155],
input_weight[156],
input_weight[157],
input_weight[158],
input_weight[159],
input_weight[160],
input_weight[161],
input_weight[162],
input_weight[163],
input_weight[164],
input_weight[165],
input_weight[166],
input_weight[167],
input_weight[168],
input_weight[169],
input_weight[170],
input_weight[171],
input_weight[172],
input_weight[173],
input_weight[174],
input_weight[175],
input_weight[176],
input_weight[177],
input_weight[178],
input_weight[179],
input_weight[180],
input_weight[181],
input_weight[182],
input_weight[183],
input_weight[184],
input_weight[185],
input_weight[186],
input_weight[187],
input_weight[188],
input_weight[189],
input_weight[190],
input_weight[191],
input_weight[192],
input_weight[193],
input_weight[194],
input_weight[195],
input_weight[196],
input_weight[197],
input_weight[198],
input_weight[199]
} = {
8'sd127,
8'sd127,
8'sd0,
8'sd127,
-8'sd128,
8'sd127,
8'sd127,
8'sd127,
-8'sd128,
8'sd127,
-8'sd128,
8'sd0,
-8'sd128,
-8'sd128,
8'sd127,
8'sd0,
-8'sd128,
-8'sd128,
-8'sd128,
-8'sd128,
8'sd0,
8'sd127,
8'sd127,
8'sd127,
8'sd127,
8'sd127,
8'sd127,
-8'sd128,
8'sd127,
-8'sd128,
8'sd127,
-8'sd128,
8'sd127,
8'sd0,
8'sd127,
8'sd127,
8'sd127,
-8'sd128,
-8'sd128,
-8'sd128,
8'sd0,
8'sd127,
8'sd127,
8'sd127,
-8'sd128,
-8'sd128,
-8'sd128,
-8'sd128,
8'sd0,
8'sd127,
8'sd127,
-8'sd128,
-8'sd128,
8'sd127,
-8'sd128,
-8'sd128,
-8'sd128,
-8'sd128,
-8'sd128,
8'sd0,
-8'sd128,
-8'sd128,
-8'sd128,
8'sd127,
-8'sd128,
-8'sd128,
8'sd127,
8'sd127,
8'sd127,
8'sd127,
-8'sd128,
8'sd127,
-8'sd128,
-8'sd128,
-8'sd128,
8'sd127,
8'sd127,
-8'sd128,
-8'sd128,
-8'sd128,
8'sd127,
-8'sd128,
-8'sd128,
-8'sd128,
-8'sd128,
-8'sd128,
8'sd0,
8'sd127,
8'sd127,
8'sd127,
8'sd127,
-8'sd128,
8'sd127,
-8'sd128,
-8'sd128,
8'sd0,
8'sd127,
-8'sd128,
8'sd127,
8'sd127,
8'sd127,
8'sd0,
-8'sd128,
8'sd0,
8'sd127,
8'sd127,
8'sd127,
-8'sd128,
8'sd0,
-8'sd128,
8'sd127,
8'sd127,
8'sd127,
-8'sd128,
8'sd127,
8'sd127,
-8'sd128,
-8'sd128,
8'sd127,
-8'sd128,
8'sd127,
-8'sd128,
-8'sd128,
8'sd127,
8'sd127,
-8'sd128,
-8'sd128,
8'sd127,
-8'sd128,
-8'sd128,
-8'sd128,
-8'sd128,
-8'sd128,
8'sd127,
8'sd127,
-8'sd128,
-8'sd128,
8'sd127,
8'sd0,
-8'sd128,
-8'sd128,
8'sd127,
8'sd127,
8'sd127,
8'sd127,
-8'sd128,
-8'sd128,
8'sd127,
8'sd127,
8'sd127,
-8'sd128,
8'sd127,
-8'sd128,
8'sd0,
8'sd127,
-8'sd128,
8'sd127,
-8'sd128,
-8'sd128,
-8'sd128,
-8'sd128,
8'sd127,
8'sd0,
-8'sd128,
8'sd0,
-8'sd128,
-8'sd128,
8'sd127,
-8'sd128,
8'sd127,
8'sd127,
-8'sd128,
8'sd127,
-8'sd128,
-8'sd128,
8'sd0,
8'sd0,
8'sd127,
8'sd127,
-8'sd128,
8'sd127,
8'sd127,
8'sd127,
8'sd0,
-8'sd128,
8'sd127,
-8'sd128,
-8'sd128,
-8'sd128,
-8'sd128,
8'sd127,
8'sd127,
8'sd127,
8'sd127,
-8'sd128,
-8'sd128,
-8'sd128,
-8'sd128,
-8'sd128,
8'sd127
};

    // Reservoir layer
    reg signed [15:0] a_scaled = 16'd-16384;
reg signed [15:0] b_scaled = 16'd16384;
reg signed [15:0] c_scaled = 16'd-19248;
reg signed [15:0] d_scaled = 16'd19248;
reg signed [31:0] reservoir_state [0: num_reservoir_neurons-1];
initial {
reservoir_state[0],
reservoir_state[1],
reservoir_state[2],
reservoir_state[3],
reservoir_state[4],
reservoir_state[5],
reservoir_state[6],
reservoir_state[7],
reservoir_state[8],
reservoir_state[9],
reservoir_state[10],
reservoir_state[11],
reservoir_state[12],
reservoir_state[13],
reservoir_state[14],
reservoir_state[15],
reservoir_state[16],
reservoir_state[17],
reservoir_state[18],
reservoir_state[19],
reservoir_state[20],
reservoir_state[21],
reservoir_state[22],
reservoir_state[23],
reservoir_state[24],
reservoir_state[25],
reservoir_state[26],
reservoir_state[27],
reservoir_state[28],
reservoir_state[29],
reservoir_state[30],
reservoir_state[31],
reservoir_state[32],
reservoir_state[33],
reservoir_state[34],
reservoir_state[35],
reservoir_state[36],
reservoir_state[37],
reservoir_state[38],
reservoir_state[39],
reservoir_state[40],
reservoir_state[41],
reservoir_state[42],
reservoir_state[43],
reservoir_state[44],
reservoir_state[45],
reservoir_state[46],
reservoir_state[47],
reservoir_state[48],
reservoir_state[49],
reservoir_state[50],
reservoir_state[51],
reservoir_state[52],
reservoir_state[53],
reservoir_state[54],
reservoir_state[55],
reservoir_state[56],
reservoir_state[57],
reservoir_state[58],
reservoir_state[59],
reservoir_state[60],
reservoir_state[61],
reservoir_state[62],
reservoir_state[63],
reservoir_state[64],
reservoir_state[65],
reservoir_state[66],
reservoir_state[67],
reservoir_state[68],
reservoir_state[69],
reservoir_state[70],
reservoir_state[71],
reservoir_state[72],
reservoir_state[73],
reservoir_state[74],
reservoir_state[75],
reservoir_state[76],
reservoir_state[77],
reservoir_state[78],
reservoir_state[79],
reservoir_state[80],
reservoir_state[81],
reservoir_state[82],
reservoir_state[83],
reservoir_state[84],
reservoir_state[85],
reservoir_state[86],
reservoir_state[87],
reservoir_state[88],
reservoir_state[89],
reservoir_state[90],
reservoir_state[91],
reservoir_state[92],
reservoir_state[93],
reservoir_state[94],
reservoir_state[95],
reservoir_state[96],
reservoir_state[97],
reservoir_state[98],
reservoir_state[99],
reservoir_state[100],
reservoir_state[101],
reservoir_state[102],
reservoir_state[103],
reservoir_state[104],
reservoir_state[105],
reservoir_state[106],
reservoir_state[107],
reservoir_state[108],
reservoir_state[109],
reservoir_state[110],
reservoir_state[111],
reservoir_state[112],
reservoir_state[113],
reservoir_state[114],
reservoir_state[115],
reservoir_state[116],
reservoir_state[117],
reservoir_state[118],
reservoir_state[119],
reservoir_state[120],
reservoir_state[121],
reservoir_state[122],
reservoir_state[123],
reservoir_state[124],
reservoir_state[125],
reservoir_state[126],
reservoir_state[127],
reservoir_state[128],
reservoir_state[129],
reservoir_state[130],
reservoir_state[131],
reservoir_state[132],
reservoir_state[133],
reservoir_state[134],
reservoir_state[135],
reservoir_state[136],
reservoir_state[137],
reservoir_state[138],
reservoir_state[139],
reservoir_state[140],
reservoir_state[141],
reservoir_state[142],
reservoir_state[143],
reservoir_state[144],
reservoir_state[145],
reservoir_state[146],
reservoir_state[147],
reservoir_state[148],
reservoir_state[149],
reservoir_state[150],
reservoir_state[151],
reservoir_state[152],
reservoir_state[153],
reservoir_state[154],
reservoir_state[155],
reservoir_state[156],
reservoir_state[157],
reservoir_state[158],
reservoir_state[159],
reservoir_state[160],
reservoir_state[161],
reservoir_state[162],
reservoir_state[163],
reservoir_state[164],
reservoir_state[165],
reservoir_state[166],
reservoir_state[167],
reservoir_state[168],
reservoir_state[169],
reservoir_state[170],
reservoir_state[171],
reservoir_state[172],
reservoir_state[173],
reservoir_state[174],
reservoir_state[175],
reservoir_state[176],
reservoir_state[177],
reservoir_state[178],
reservoir_state[179],
reservoir_state[180],
reservoir_state[181],
reservoir_state[182],
reservoir_state[183],
reservoir_state[184],
reservoir_state[185],
reservoir_state[186],
reservoir_state[187],
reservoir_state[188],
reservoir_state[189],
reservoir_state[190],
reservoir_state[191],
reservoir_state[192],
reservoir_state[193],
reservoir_state[194],
reservoir_state[195],
reservoir_state[196],
reservoir_state[197],
reservoir_state[198],
reservoir_state[199]
} = {
-32'sd84,
-32'sd80,
-32'sd124,
-32'sd55,
32'sd121,
32'sd112,
32'sd94,
32'sd115,
32'sd116,
-32'sd115,
32'sd101,
-32'sd58,
-32'sd77,
-32'sd119,
-32'sd101,
32'sd61,
32'sd71,
32'sd54,
32'sd116,
-32'sd95,
-32'sd101,
-32'sd122,
-32'sd113,
-32'sd101,
-32'sd121,
32'sd31,
32'sd124,
-32'sd5,
-32'sd126,
32'sd101,
32'sd70,
-32'sd6,
-32'sd94,
32'sd124,
32'sd84,
-32'sd124,
32'sd105,
-32'sd69,
32'sd89,
-32'sd33,
-32'sd65,
32'sd109,
-32'sd126,
32'sd76,
32'sd81,
32'sd111,
-32'sd84,
32'sd62,
32'sd111,
-32'sd105,
32'sd120,
32'sd115,
32'sd90,
32'sd38,
32'sd127,
-32'sd126,
-32'sd43,
-32'sd86,
32'sd122,
-32'sd29,
-32'sd110,
32'sd14,
-32'sd89,
-32'sd107,
32'sd1,
32'sd117,
32'sd124,
32'sd108,
32'sd115,
32'sd108,
-32'sd82,
32'sd60,
-32'sd40,
-32'sd118,
32'sd72,
-32'sd107,
32'sd67,
32'sd117,
-32'sd121,
32'sd104,
32'sd77,
32'sd119,
32'sd112,
32'sd83,
-32'sd125,
32'sd92,
32'sd9,
32'sd91,
32'sd114,
-32'sd123,
-32'sd90,
-32'sd9,
32'sd127,
-32'sd77,
32'sd105,
32'sd46,
-32'sd62,
-32'sd106,
32'sd87,
-32'sd104,
-32'sd82,
-32'sd88,
32'sd126,
-32'sd64,
32'sd11,
32'sd116,
-32'sd126,
32'sd87,
32'sd96,
32'sd80,
-32'sd116,
-32'sd80,
32'sd119,
32'sd115,
-32'sd45,
32'sd38,
-32'sd24,
-32'sd111,
32'sd114,
-32'sd111,
32'sd103,
32'sd51,
-32'sd82,
32'sd58,
32'sd23,
-32'sd61,
-32'sd119,
32'sd10,
-32'sd117,
32'sd112,
-32'sd34,
-32'sd100,
32'sd82,
32'sd127,
32'sd32,
32'sd93,
-32'sd110,
32'sd79,
-32'sd20,
32'sd52,
-32'sd71,
-32'sd124,
-32'sd10,
32'sd119,
-32'sd105,
32'sd14,
32'sd122,
-32'sd46,
-32'sd121,
32'sd100,
32'sd71,
-32'sd99,
32'sd104,
32'sd73,
-32'sd104,
-32'sd127,
-32'sd111,
-32'sd93,
32'sd26,
-32'sd87,
-32'sd7,
-32'sd92,
32'sd89,
-32'sd16,
-32'sd43,
-32'sd107,
-32'sd122,
32'sd127,
32'sd111,
-32'sd123,
32'sd8,
32'sd126,
-32'sd123,
32'sd16,
-32'sd127,
-32'sd116,
32'sd65,
32'sd126,
32'sd112,
32'sd118,
32'sd71,
-32'sd106,
32'sd23,
32'sd60,
32'sd127,
32'sd104,
32'sd107,
-32'sd85,
-32'sd108,
-32'sd68,
-32'sd82,
32'sd98,
32'sd114,
32'sd119,
32'sd110,
32'sd57,
-32'sd78,
32'sd19,
-32'sd128,
-32'sd92
};reg signed [7:0] reservoir_weight [0: num_reservoir_neurons-1][0: num_reservoir_neurons-1];initial {
{reservoir_weight[0][0],
reservoir_weight[0][1],
reservoir_weight[0][2],
reservoir_weight[0][3],
reservoir_weight[0][4],
reservoir_weight[0][5],
reservoir_weight[0][6],
reservoir_weight[0][7],
reservoir_weight[0][8],
reservoir_weight[0][9],
reservoir_weight[0][10],
reservoir_weight[0][11],
reservoir_weight[0][12],
reservoir_weight[0][13],
reservoir_weight[0][14],
reservoir_weight[0][15],
reservoir_weight[0][16],
reservoir_weight[0][17],
reservoir_weight[0][18],
reservoir_weight[0][19],
reservoir_weight[0][20],
reservoir_weight[0][21],
reservoir_weight[0][22],
reservoir_weight[0][23],
reservoir_weight[0][24],
reservoir_weight[0][25],
reservoir_weight[0][26],
reservoir_weight[0][27],
reservoir_weight[0][28],
reservoir_weight[0][29],
reservoir_weight[0][30],
reservoir_weight[0][31],
reservoir_weight[0][32],
reservoir_weight[0][33],
reservoir_weight[0][34],
reservoir_weight[0][35],
reservoir_weight[0][36],
reservoir_weight[0][37],
reservoir_weight[0][38],
reservoir_weight[0][39],
reservoir_weight[0][40],
reservoir_weight[0][41],
reservoir_weight[0][42],
reservoir_weight[0][43],
reservoir_weight[0][44],
reservoir_weight[0][45],
reservoir_weight[0][46],
reservoir_weight[0][47],
reservoir_weight[0][48],
reservoir_weight[0][49],
reservoir_weight[0][50],
reservoir_weight[0][51],
reservoir_weight[0][52],
reservoir_weight[0][53],
reservoir_weight[0][54],
reservoir_weight[0][55],
reservoir_weight[0][56],
reservoir_weight[0][57],
reservoir_weight[0][58],
reservoir_weight[0][59],
reservoir_weight[0][60],
reservoir_weight[0][61],
reservoir_weight[0][62],
reservoir_weight[0][63],
reservoir_weight[0][64],
reservoir_weight[0][65],
reservoir_weight[0][66],
reservoir_weight[0][67],
reservoir_weight[0][68],
reservoir_weight[0][69],
reservoir_weight[0][70],
reservoir_weight[0][71],
reservoir_weight[0][72],
reservoir_weight[0][73],
reservoir_weight[0][74],
reservoir_weight[0][75],
reservoir_weight[0][76],
reservoir_weight[0][77],
reservoir_weight[0][78],
reservoir_weight[0][79],
reservoir_weight[0][80],
reservoir_weight[0][81],
reservoir_weight[0][82],
reservoir_weight[0][83],
reservoir_weight[0][84],
reservoir_weight[0][85],
reservoir_weight[0][86],
reservoir_weight[0][87],
reservoir_weight[0][88],
reservoir_weight[0][89],
reservoir_weight[0][90],
reservoir_weight[0][91],
reservoir_weight[0][92],
reservoir_weight[0][93],
reservoir_weight[0][94],
reservoir_weight[0][95],
reservoir_weight[0][96],
reservoir_weight[0][97],
reservoir_weight[0][98],
reservoir_weight[0][99],
reservoir_weight[0][100],
reservoir_weight[0][101],
reservoir_weight[0][102],
reservoir_weight[0][103],
reservoir_weight[0][104],
reservoir_weight[0][105],
reservoir_weight[0][106],
reservoir_weight[0][107],
reservoir_weight[0][108],
reservoir_weight[0][109],
reservoir_weight[0][110],
reservoir_weight[0][111],
reservoir_weight[0][112],
reservoir_weight[0][113],
reservoir_weight[0][114],
reservoir_weight[0][115],
reservoir_weight[0][116],
reservoir_weight[0][117],
reservoir_weight[0][118],
reservoir_weight[0][119],
reservoir_weight[0][120],
reservoir_weight[0][121],
reservoir_weight[0][122],
reservoir_weight[0][123],
reservoir_weight[0][124],
reservoir_weight[0][125],
reservoir_weight[0][126],
reservoir_weight[0][127],
reservoir_weight[0][128],
reservoir_weight[0][129],
reservoir_weight[0][130],
reservoir_weight[0][131],
reservoir_weight[0][132],
reservoir_weight[0][133],
reservoir_weight[0][134],
reservoir_weight[0][135],
reservoir_weight[0][136],
reservoir_weight[0][137],
reservoir_weight[0][138],
reservoir_weight[0][139],
reservoir_weight[0][140],
reservoir_weight[0][141],
reservoir_weight[0][142],
reservoir_weight[0][143],
reservoir_weight[0][144],
reservoir_weight[0][145],
reservoir_weight[0][146],
reservoir_weight[0][147],
reservoir_weight[0][148],
reservoir_weight[0][149],
reservoir_weight[0][150],
reservoir_weight[0][151],
reservoir_weight[0][152],
reservoir_weight[0][153],
reservoir_weight[0][154],
reservoir_weight[0][155],
reservoir_weight[0][156],
reservoir_weight[0][157],
reservoir_weight[0][158],
reservoir_weight[0][159],
reservoir_weight[0][160],
reservoir_weight[0][161],
reservoir_weight[0][162],
reservoir_weight[0][163],
reservoir_weight[0][164],
reservoir_weight[0][165],
reservoir_weight[0][166],
reservoir_weight[0][167],
reservoir_weight[0][168],
reservoir_weight[0][169],
reservoir_weight[0][170],
reservoir_weight[0][171],
reservoir_weight[0][172],
reservoir_weight[0][173],
reservoir_weight[0][174],
reservoir_weight[0][175],
reservoir_weight[0][176],
reservoir_weight[0][177],
reservoir_weight[0][178],
reservoir_weight[0][179],
reservoir_weight[0][180],
reservoir_weight[0][181],
reservoir_weight[0][182],
reservoir_weight[0][183],
reservoir_weight[0][184],
reservoir_weight[0][185],
reservoir_weight[0][186],
reservoir_weight[0][187],
reservoir_weight[0][188],
reservoir_weight[0][189],
reservoir_weight[0][190],
reservoir_weight[0][191],
reservoir_weight[0][192],
reservoir_weight[0][193],
reservoir_weight[0][194],
reservoir_weight[0][195],
reservoir_weight[0][196],
reservoir_weight[0][197],
reservoir_weight[0][198],
reservoir_weight[0][199]
},
{reservoir_weight[1][0],
reservoir_weight[1][1],
reservoir_weight[1][2],
reservoir_weight[1][3],
reservoir_weight[1][4],
reservoir_weight[1][5],
reservoir_weight[1][6],
reservoir_weight[1][7],
reservoir_weight[1][8],
reservoir_weight[1][9],
reservoir_weight[1][10],
reservoir_weight[1][11],
reservoir_weight[1][12],
reservoir_weight[1][13],
reservoir_weight[1][14],
reservoir_weight[1][15],
reservoir_weight[1][16],
reservoir_weight[1][17],
reservoir_weight[1][18],
reservoir_weight[1][19],
reservoir_weight[1][20],
reservoir_weight[1][21],
reservoir_weight[1][22],
reservoir_weight[1][23],
reservoir_weight[1][24],
reservoir_weight[1][25],
reservoir_weight[1][26],
reservoir_weight[1][27],
reservoir_weight[1][28],
reservoir_weight[1][29],
reservoir_weight[1][30],
reservoir_weight[1][31],
reservoir_weight[1][32],
reservoir_weight[1][33],
reservoir_weight[1][34],
reservoir_weight[1][35],
reservoir_weight[1][36],
reservoir_weight[1][37],
reservoir_weight[1][38],
reservoir_weight[1][39],
reservoir_weight[1][40],
reservoir_weight[1][41],
reservoir_weight[1][42],
reservoir_weight[1][43],
reservoir_weight[1][44],
reservoir_weight[1][45],
reservoir_weight[1][46],
reservoir_weight[1][47],
reservoir_weight[1][48],
reservoir_weight[1][49],
reservoir_weight[1][50],
reservoir_weight[1][51],
reservoir_weight[1][52],
reservoir_weight[1][53],
reservoir_weight[1][54],
reservoir_weight[1][55],
reservoir_weight[1][56],
reservoir_weight[1][57],
reservoir_weight[1][58],
reservoir_weight[1][59],
reservoir_weight[1][60],
reservoir_weight[1][61],
reservoir_weight[1][62],
reservoir_weight[1][63],
reservoir_weight[1][64],
reservoir_weight[1][65],
reservoir_weight[1][66],
reservoir_weight[1][67],
reservoir_weight[1][68],
reservoir_weight[1][69],
reservoir_weight[1][70],
reservoir_weight[1][71],
reservoir_weight[1][72],
reservoir_weight[1][73],
reservoir_weight[1][74],
reservoir_weight[1][75],
reservoir_weight[1][76],
reservoir_weight[1][77],
reservoir_weight[1][78],
reservoir_weight[1][79],
reservoir_weight[1][80],
reservoir_weight[1][81],
reservoir_weight[1][82],
reservoir_weight[1][83],
reservoir_weight[1][84],
reservoir_weight[1][85],
reservoir_weight[1][86],
reservoir_weight[1][87],
reservoir_weight[1][88],
reservoir_weight[1][89],
reservoir_weight[1][90],
reservoir_weight[1][91],
reservoir_weight[1][92],
reservoir_weight[1][93],
reservoir_weight[1][94],
reservoir_weight[1][95],
reservoir_weight[1][96],
reservoir_weight[1][97],
reservoir_weight[1][98],
reservoir_weight[1][99],
reservoir_weight[1][100],
reservoir_weight[1][101],
reservoir_weight[1][102],
reservoir_weight[1][103],
reservoir_weight[1][104],
reservoir_weight[1][105],
reservoir_weight[1][106],
reservoir_weight[1][107],
reservoir_weight[1][108],
reservoir_weight[1][109],
reservoir_weight[1][110],
reservoir_weight[1][111],
reservoir_weight[1][112],
reservoir_weight[1][113],
reservoir_weight[1][114],
reservoir_weight[1][115],
reservoir_weight[1][116],
reservoir_weight[1][117],
reservoir_weight[1][118],
reservoir_weight[1][119],
reservoir_weight[1][120],
reservoir_weight[1][121],
reservoir_weight[1][122],
reservoir_weight[1][123],
reservoir_weight[1][124],
reservoir_weight[1][125],
reservoir_weight[1][126],
reservoir_weight[1][127],
reservoir_weight[1][128],
reservoir_weight[1][129],
reservoir_weight[1][130],
reservoir_weight[1][131],
reservoir_weight[1][132],
reservoir_weight[1][133],
reservoir_weight[1][134],
reservoir_weight[1][135],
reservoir_weight[1][136],
reservoir_weight[1][137],
reservoir_weight[1][138],
reservoir_weight[1][139],
reservoir_weight[1][140],
reservoir_weight[1][141],
reservoir_weight[1][142],
reservoir_weight[1][143],
reservoir_weight[1][144],
reservoir_weight[1][145],
reservoir_weight[1][146],
reservoir_weight[1][147],
reservoir_weight[1][148],
reservoir_weight[1][149],
reservoir_weight[1][150],
reservoir_weight[1][151],
reservoir_weight[1][152],
reservoir_weight[1][153],
reservoir_weight[1][154],
reservoir_weight[1][155],
reservoir_weight[1][156],
reservoir_weight[1][157],
reservoir_weight[1][158],
reservoir_weight[1][159],
reservoir_weight[1][160],
reservoir_weight[1][161],
reservoir_weight[1][162],
reservoir_weight[1][163],
reservoir_weight[1][164],
reservoir_weight[1][165],
reservoir_weight[1][166],
reservoir_weight[1][167],
reservoir_weight[1][168],
reservoir_weight[1][169],
reservoir_weight[1][170],
reservoir_weight[1][171],
reservoir_weight[1][172],
reservoir_weight[1][173],
reservoir_weight[1][174],
reservoir_weight[1][175],
reservoir_weight[1][176],
reservoir_weight[1][177],
reservoir_weight[1][178],
reservoir_weight[1][179],
reservoir_weight[1][180],
reservoir_weight[1][181],
reservoir_weight[1][182],
reservoir_weight[1][183],
reservoir_weight[1][184],
reservoir_weight[1][185],
reservoir_weight[1][186],
reservoir_weight[1][187],
reservoir_weight[1][188],
reservoir_weight[1][189],
reservoir_weight[1][190],
reservoir_weight[1][191],
reservoir_weight[1][192],
reservoir_weight[1][193],
reservoir_weight[1][194],
reservoir_weight[1][195],
reservoir_weight[1][196],
reservoir_weight[1][197],
reservoir_weight[1][198],
reservoir_weight[1][199]
},
{reservoir_weight[2][0],
reservoir_weight[2][1],
reservoir_weight[2][2],
reservoir_weight[2][3],
reservoir_weight[2][4],
reservoir_weight[2][5],
reservoir_weight[2][6],
reservoir_weight[2][7],
reservoir_weight[2][8],
reservoir_weight[2][9],
reservoir_weight[2][10],
reservoir_weight[2][11],
reservoir_weight[2][12],
reservoir_weight[2][13],
reservoir_weight[2][14],
reservoir_weight[2][15],
reservoir_weight[2][16],
reservoir_weight[2][17],
reservoir_weight[2][18],
reservoir_weight[2][19],
reservoir_weight[2][20],
reservoir_weight[2][21],
reservoir_weight[2][22],
reservoir_weight[2][23],
reservoir_weight[2][24],
reservoir_weight[2][25],
reservoir_weight[2][26],
reservoir_weight[2][27],
reservoir_weight[2][28],
reservoir_weight[2][29],
reservoir_weight[2][30],
reservoir_weight[2][31],
reservoir_weight[2][32],
reservoir_weight[2][33],
reservoir_weight[2][34],
reservoir_weight[2][35],
reservoir_weight[2][36],
reservoir_weight[2][37],
reservoir_weight[2][38],
reservoir_weight[2][39],
reservoir_weight[2][40],
reservoir_weight[2][41],
reservoir_weight[2][42],
reservoir_weight[2][43],
reservoir_weight[2][44],
reservoir_weight[2][45],
reservoir_weight[2][46],
reservoir_weight[2][47],
reservoir_weight[2][48],
reservoir_weight[2][49],
reservoir_weight[2][50],
reservoir_weight[2][51],
reservoir_weight[2][52],
reservoir_weight[2][53],
reservoir_weight[2][54],
reservoir_weight[2][55],
reservoir_weight[2][56],
reservoir_weight[2][57],
reservoir_weight[2][58],
reservoir_weight[2][59],
reservoir_weight[2][60],
reservoir_weight[2][61],
reservoir_weight[2][62],
reservoir_weight[2][63],
reservoir_weight[2][64],
reservoir_weight[2][65],
reservoir_weight[2][66],
reservoir_weight[2][67],
reservoir_weight[2][68],
reservoir_weight[2][69],
reservoir_weight[2][70],
reservoir_weight[2][71],
reservoir_weight[2][72],
reservoir_weight[2][73],
reservoir_weight[2][74],
reservoir_weight[2][75],
reservoir_weight[2][76],
reservoir_weight[2][77],
reservoir_weight[2][78],
reservoir_weight[2][79],
reservoir_weight[2][80],
reservoir_weight[2][81],
reservoir_weight[2][82],
reservoir_weight[2][83],
reservoir_weight[2][84],
reservoir_weight[2][85],
reservoir_weight[2][86],
reservoir_weight[2][87],
reservoir_weight[2][88],
reservoir_weight[2][89],
reservoir_weight[2][90],
reservoir_weight[2][91],
reservoir_weight[2][92],
reservoir_weight[2][93],
reservoir_weight[2][94],
reservoir_weight[2][95],
reservoir_weight[2][96],
reservoir_weight[2][97],
reservoir_weight[2][98],
reservoir_weight[2][99],
reservoir_weight[2][100],
reservoir_weight[2][101],
reservoir_weight[2][102],
reservoir_weight[2][103],
reservoir_weight[2][104],
reservoir_weight[2][105],
reservoir_weight[2][106],
reservoir_weight[2][107],
reservoir_weight[2][108],
reservoir_weight[2][109],
reservoir_weight[2][110],
reservoir_weight[2][111],
reservoir_weight[2][112],
reservoir_weight[2][113],
reservoir_weight[2][114],
reservoir_weight[2][115],
reservoir_weight[2][116],
reservoir_weight[2][117],
reservoir_weight[2][118],
reservoir_weight[2][119],
reservoir_weight[2][120],
reservoir_weight[2][121],
reservoir_weight[2][122],
reservoir_weight[2][123],
reservoir_weight[2][124],
reservoir_weight[2][125],
reservoir_weight[2][126],
reservoir_weight[2][127],
reservoir_weight[2][128],
reservoir_weight[2][129],
reservoir_weight[2][130],
reservoir_weight[2][131],
reservoir_weight[2][132],
reservoir_weight[2][133],
reservoir_weight[2][134],
reservoir_weight[2][135],
reservoir_weight[2][136],
reservoir_weight[2][137],
reservoir_weight[2][138],
reservoir_weight[2][139],
reservoir_weight[2][140],
reservoir_weight[2][141],
reservoir_weight[2][142],
reservoir_weight[2][143],
reservoir_weight[2][144],
reservoir_weight[2][145],
reservoir_weight[2][146],
reservoir_weight[2][147],
reservoir_weight[2][148],
reservoir_weight[2][149],
reservoir_weight[2][150],
reservoir_weight[2][151],
reservoir_weight[2][152],
reservoir_weight[2][153],
reservoir_weight[2][154],
reservoir_weight[2][155],
reservoir_weight[2][156],
reservoir_weight[2][157],
reservoir_weight[2][158],
reservoir_weight[2][159],
reservoir_weight[2][160],
reservoir_weight[2][161],
reservoir_weight[2][162],
reservoir_weight[2][163],
reservoir_weight[2][164],
reservoir_weight[2][165],
reservoir_weight[2][166],
reservoir_weight[2][167],
reservoir_weight[2][168],
reservoir_weight[2][169],
reservoir_weight[2][170],
reservoir_weight[2][171],
reservoir_weight[2][172],
reservoir_weight[2][173],
reservoir_weight[2][174],
reservoir_weight[2][175],
reservoir_weight[2][176],
reservoir_weight[2][177],
reservoir_weight[2][178],
reservoir_weight[2][179],
reservoir_weight[2][180],
reservoir_weight[2][181],
reservoir_weight[2][182],
reservoir_weight[2][183],
reservoir_weight[2][184],
reservoir_weight[2][185],
reservoir_weight[2][186],
reservoir_weight[2][187],
reservoir_weight[2][188],
reservoir_weight[2][189],
reservoir_weight[2][190],
reservoir_weight[2][191],
reservoir_weight[2][192],
reservoir_weight[2][193],
reservoir_weight[2][194],
reservoir_weight[2][195],
reservoir_weight[2][196],
reservoir_weight[2][197],
reservoir_weight[2][198],
reservoir_weight[2][199]
},
{reservoir_weight[3][0],
reservoir_weight[3][1],
reservoir_weight[3][2],
reservoir_weight[3][3],
reservoir_weight[3][4],
reservoir_weight[3][5],
reservoir_weight[3][6],
reservoir_weight[3][7],
reservoir_weight[3][8],
reservoir_weight[3][9],
reservoir_weight[3][10],
reservoir_weight[3][11],
reservoir_weight[3][12],
reservoir_weight[3][13],
reservoir_weight[3][14],
reservoir_weight[3][15],
reservoir_weight[3][16],
reservoir_weight[3][17],
reservoir_weight[3][18],
reservoir_weight[3][19],
reservoir_weight[3][20],
reservoir_weight[3][21],
reservoir_weight[3][22],
reservoir_weight[3][23],
reservoir_weight[3][24],
reservoir_weight[3][25],
reservoir_weight[3][26],
reservoir_weight[3][27],
reservoir_weight[3][28],
reservoir_weight[3][29],
reservoir_weight[3][30],
reservoir_weight[3][31],
reservoir_weight[3][32],
reservoir_weight[3][33],
reservoir_weight[3][34],
reservoir_weight[3][35],
reservoir_weight[3][36],
reservoir_weight[3][37],
reservoir_weight[3][38],
reservoir_weight[3][39],
reservoir_weight[3][40],
reservoir_weight[3][41],
reservoir_weight[3][42],
reservoir_weight[3][43],
reservoir_weight[3][44],
reservoir_weight[3][45],
reservoir_weight[3][46],
reservoir_weight[3][47],
reservoir_weight[3][48],
reservoir_weight[3][49],
reservoir_weight[3][50],
reservoir_weight[3][51],
reservoir_weight[3][52],
reservoir_weight[3][53],
reservoir_weight[3][54],
reservoir_weight[3][55],
reservoir_weight[3][56],
reservoir_weight[3][57],
reservoir_weight[3][58],
reservoir_weight[3][59],
reservoir_weight[3][60],
reservoir_weight[3][61],
reservoir_weight[3][62],
reservoir_weight[3][63],
reservoir_weight[3][64],
reservoir_weight[3][65],
reservoir_weight[3][66],
reservoir_weight[3][67],
reservoir_weight[3][68],
reservoir_weight[3][69],
reservoir_weight[3][70],
reservoir_weight[3][71],
reservoir_weight[3][72],
reservoir_weight[3][73],
reservoir_weight[3][74],
reservoir_weight[3][75],
reservoir_weight[3][76],
reservoir_weight[3][77],
reservoir_weight[3][78],
reservoir_weight[3][79],
reservoir_weight[3][80],
reservoir_weight[3][81],
reservoir_weight[3][82],
reservoir_weight[3][83],
reservoir_weight[3][84],
reservoir_weight[3][85],
reservoir_weight[3][86],
reservoir_weight[3][87],
reservoir_weight[3][88],
reservoir_weight[3][89],
reservoir_weight[3][90],
reservoir_weight[3][91],
reservoir_weight[3][92],
reservoir_weight[3][93],
reservoir_weight[3][94],
reservoir_weight[3][95],
reservoir_weight[3][96],
reservoir_weight[3][97],
reservoir_weight[3][98],
reservoir_weight[3][99],
reservoir_weight[3][100],
reservoir_weight[3][101],
reservoir_weight[3][102],
reservoir_weight[3][103],
reservoir_weight[3][104],
reservoir_weight[3][105],
reservoir_weight[3][106],
reservoir_weight[3][107],
reservoir_weight[3][108],
reservoir_weight[3][109],
reservoir_weight[3][110],
reservoir_weight[3][111],
reservoir_weight[3][112],
reservoir_weight[3][113],
reservoir_weight[3][114],
reservoir_weight[3][115],
reservoir_weight[3][116],
reservoir_weight[3][117],
reservoir_weight[3][118],
reservoir_weight[3][119],
reservoir_weight[3][120],
reservoir_weight[3][121],
reservoir_weight[3][122],
reservoir_weight[3][123],
reservoir_weight[3][124],
reservoir_weight[3][125],
reservoir_weight[3][126],
reservoir_weight[3][127],
reservoir_weight[3][128],
reservoir_weight[3][129],
reservoir_weight[3][130],
reservoir_weight[3][131],
reservoir_weight[3][132],
reservoir_weight[3][133],
reservoir_weight[3][134],
reservoir_weight[3][135],
reservoir_weight[3][136],
reservoir_weight[3][137],
reservoir_weight[3][138],
reservoir_weight[3][139],
reservoir_weight[3][140],
reservoir_weight[3][141],
reservoir_weight[3][142],
reservoir_weight[3][143],
reservoir_weight[3][144],
reservoir_weight[3][145],
reservoir_weight[3][146],
reservoir_weight[3][147],
reservoir_weight[3][148],
reservoir_weight[3][149],
reservoir_weight[3][150],
reservoir_weight[3][151],
reservoir_weight[3][152],
reservoir_weight[3][153],
reservoir_weight[3][154],
reservoir_weight[3][155],
reservoir_weight[3][156],
reservoir_weight[3][157],
reservoir_weight[3][158],
reservoir_weight[3][159],
reservoir_weight[3][160],
reservoir_weight[3][161],
reservoir_weight[3][162],
reservoir_weight[3][163],
reservoir_weight[3][164],
reservoir_weight[3][165],
reservoir_weight[3][166],
reservoir_weight[3][167],
reservoir_weight[3][168],
reservoir_weight[3][169],
reservoir_weight[3][170],
reservoir_weight[3][171],
reservoir_weight[3][172],
reservoir_weight[3][173],
reservoir_weight[3][174],
reservoir_weight[3][175],
reservoir_weight[3][176],
reservoir_weight[3][177],
reservoir_weight[3][178],
reservoir_weight[3][179],
reservoir_weight[3][180],
reservoir_weight[3][181],
reservoir_weight[3][182],
reservoir_weight[3][183],
reservoir_weight[3][184],
reservoir_weight[3][185],
reservoir_weight[3][186],
reservoir_weight[3][187],
reservoir_weight[3][188],
reservoir_weight[3][189],
reservoir_weight[3][190],
reservoir_weight[3][191],
reservoir_weight[3][192],
reservoir_weight[3][193],
reservoir_weight[3][194],
reservoir_weight[3][195],
reservoir_weight[3][196],
reservoir_weight[3][197],
reservoir_weight[3][198],
reservoir_weight[3][199]
},
{reservoir_weight[4][0],
reservoir_weight[4][1],
reservoir_weight[4][2],
reservoir_weight[4][3],
reservoir_weight[4][4],
reservoir_weight[4][5],
reservoir_weight[4][6],
reservoir_weight[4][7],
reservoir_weight[4][8],
reservoir_weight[4][9],
reservoir_weight[4][10],
reservoir_weight[4][11],
reservoir_weight[4][12],
reservoir_weight[4][13],
reservoir_weight[4][14],
reservoir_weight[4][15],
reservoir_weight[4][16],
reservoir_weight[4][17],
reservoir_weight[4][18],
reservoir_weight[4][19],
reservoir_weight[4][20],
reservoir_weight[4][21],
reservoir_weight[4][22],
reservoir_weight[4][23],
reservoir_weight[4][24],
reservoir_weight[4][25],
reservoir_weight[4][26],
reservoir_weight[4][27],
reservoir_weight[4][28],
reservoir_weight[4][29],
reservoir_weight[4][30],
reservoir_weight[4][31],
reservoir_weight[4][32],
reservoir_weight[4][33],
reservoir_weight[4][34],
reservoir_weight[4][35],
reservoir_weight[4][36],
reservoir_weight[4][37],
reservoir_weight[4][38],
reservoir_weight[4][39],
reservoir_weight[4][40],
reservoir_weight[4][41],
reservoir_weight[4][42],
reservoir_weight[4][43],
reservoir_weight[4][44],
reservoir_weight[4][45],
reservoir_weight[4][46],
reservoir_weight[4][47],
reservoir_weight[4][48],
reservoir_weight[4][49],
reservoir_weight[4][50],
reservoir_weight[4][51],
reservoir_weight[4][52],
reservoir_weight[4][53],
reservoir_weight[4][54],
reservoir_weight[4][55],
reservoir_weight[4][56],
reservoir_weight[4][57],
reservoir_weight[4][58],
reservoir_weight[4][59],
reservoir_weight[4][60],
reservoir_weight[4][61],
reservoir_weight[4][62],
reservoir_weight[4][63],
reservoir_weight[4][64],
reservoir_weight[4][65],
reservoir_weight[4][66],
reservoir_weight[4][67],
reservoir_weight[4][68],
reservoir_weight[4][69],
reservoir_weight[4][70],
reservoir_weight[4][71],
reservoir_weight[4][72],
reservoir_weight[4][73],
reservoir_weight[4][74],
reservoir_weight[4][75],
reservoir_weight[4][76],
reservoir_weight[4][77],
reservoir_weight[4][78],
reservoir_weight[4][79],
reservoir_weight[4][80],
reservoir_weight[4][81],
reservoir_weight[4][82],
reservoir_weight[4][83],
reservoir_weight[4][84],
reservoir_weight[4][85],
reservoir_weight[4][86],
reservoir_weight[4][87],
reservoir_weight[4][88],
reservoir_weight[4][89],
reservoir_weight[4][90],
reservoir_weight[4][91],
reservoir_weight[4][92],
reservoir_weight[4][93],
reservoir_weight[4][94],
reservoir_weight[4][95],
reservoir_weight[4][96],
reservoir_weight[4][97],
reservoir_weight[4][98],
reservoir_weight[4][99],
reservoir_weight[4][100],
reservoir_weight[4][101],
reservoir_weight[4][102],
reservoir_weight[4][103],
reservoir_weight[4][104],
reservoir_weight[4][105],
reservoir_weight[4][106],
reservoir_weight[4][107],
reservoir_weight[4][108],
reservoir_weight[4][109],
reservoir_weight[4][110],
reservoir_weight[4][111],
reservoir_weight[4][112],
reservoir_weight[4][113],
reservoir_weight[4][114],
reservoir_weight[4][115],
reservoir_weight[4][116],
reservoir_weight[4][117],
reservoir_weight[4][118],
reservoir_weight[4][119],
reservoir_weight[4][120],
reservoir_weight[4][121],
reservoir_weight[4][122],
reservoir_weight[4][123],
reservoir_weight[4][124],
reservoir_weight[4][125],
reservoir_weight[4][126],
reservoir_weight[4][127],
reservoir_weight[4][128],
reservoir_weight[4][129],
reservoir_weight[4][130],
reservoir_weight[4][131],
reservoir_weight[4][132],
reservoir_weight[4][133],
reservoir_weight[4][134],
reservoir_weight[4][135],
reservoir_weight[4][136],
reservoir_weight[4][137],
reservoir_weight[4][138],
reservoir_weight[4][139],
reservoir_weight[4][140],
reservoir_weight[4][141],
reservoir_weight[4][142],
reservoir_weight[4][143],
reservoir_weight[4][144],
reservoir_weight[4][145],
reservoir_weight[4][146],
reservoir_weight[4][147],
reservoir_weight[4][148],
reservoir_weight[4][149],
reservoir_weight[4][150],
reservoir_weight[4][151],
reservoir_weight[4][152],
reservoir_weight[4][153],
reservoir_weight[4][154],
reservoir_weight[4][155],
reservoir_weight[4][156],
reservoir_weight[4][157],
reservoir_weight[4][158],
reservoir_weight[4][159],
reservoir_weight[4][160],
reservoir_weight[4][161],
reservoir_weight[4][162],
reservoir_weight[4][163],
reservoir_weight[4][164],
reservoir_weight[4][165],
reservoir_weight[4][166],
reservoir_weight[4][167],
reservoir_weight[4][168],
reservoir_weight[4][169],
reservoir_weight[4][170],
reservoir_weight[4][171],
reservoir_weight[4][172],
reservoir_weight[4][173],
reservoir_weight[4][174],
reservoir_weight[4][175],
reservoir_weight[4][176],
reservoir_weight[4][177],
reservoir_weight[4][178],
reservoir_weight[4][179],
reservoir_weight[4][180],
reservoir_weight[4][181],
reservoir_weight[4][182],
reservoir_weight[4][183],
reservoir_weight[4][184],
reservoir_weight[4][185],
reservoir_weight[4][186],
reservoir_weight[4][187],
reservoir_weight[4][188],
reservoir_weight[4][189],
reservoir_weight[4][190],
reservoir_weight[4][191],
reservoir_weight[4][192],
reservoir_weight[4][193],
reservoir_weight[4][194],
reservoir_weight[4][195],
reservoir_weight[4][196],
reservoir_weight[4][197],
reservoir_weight[4][198],
reservoir_weight[4][199]
},
{reservoir_weight[5][0],
reservoir_weight[5][1],
reservoir_weight[5][2],
reservoir_weight[5][3],
reservoir_weight[5][4],
reservoir_weight[5][5],
reservoir_weight[5][6],
reservoir_weight[5][7],
reservoir_weight[5][8],
reservoir_weight[5][9],
reservoir_weight[5][10],
reservoir_weight[5][11],
reservoir_weight[5][12],
reservoir_weight[5][13],
reservoir_weight[5][14],
reservoir_weight[5][15],
reservoir_weight[5][16],
reservoir_weight[5][17],
reservoir_weight[5][18],
reservoir_weight[5][19],
reservoir_weight[5][20],
reservoir_weight[5][21],
reservoir_weight[5][22],
reservoir_weight[5][23],
reservoir_weight[5][24],
reservoir_weight[5][25],
reservoir_weight[5][26],
reservoir_weight[5][27],
reservoir_weight[5][28],
reservoir_weight[5][29],
reservoir_weight[5][30],
reservoir_weight[5][31],
reservoir_weight[5][32],
reservoir_weight[5][33],
reservoir_weight[5][34],
reservoir_weight[5][35],
reservoir_weight[5][36],
reservoir_weight[5][37],
reservoir_weight[5][38],
reservoir_weight[5][39],
reservoir_weight[5][40],
reservoir_weight[5][41],
reservoir_weight[5][42],
reservoir_weight[5][43],
reservoir_weight[5][44],
reservoir_weight[5][45],
reservoir_weight[5][46],
reservoir_weight[5][47],
reservoir_weight[5][48],
reservoir_weight[5][49],
reservoir_weight[5][50],
reservoir_weight[5][51],
reservoir_weight[5][52],
reservoir_weight[5][53],
reservoir_weight[5][54],
reservoir_weight[5][55],
reservoir_weight[5][56],
reservoir_weight[5][57],
reservoir_weight[5][58],
reservoir_weight[5][59],
reservoir_weight[5][60],
reservoir_weight[5][61],
reservoir_weight[5][62],
reservoir_weight[5][63],
reservoir_weight[5][64],
reservoir_weight[5][65],
reservoir_weight[5][66],
reservoir_weight[5][67],
reservoir_weight[5][68],
reservoir_weight[5][69],
reservoir_weight[5][70],
reservoir_weight[5][71],
reservoir_weight[5][72],
reservoir_weight[5][73],
reservoir_weight[5][74],
reservoir_weight[5][75],
reservoir_weight[5][76],
reservoir_weight[5][77],
reservoir_weight[5][78],
reservoir_weight[5][79],
reservoir_weight[5][80],
reservoir_weight[5][81],
reservoir_weight[5][82],
reservoir_weight[5][83],
reservoir_weight[5][84],
reservoir_weight[5][85],
reservoir_weight[5][86],
reservoir_weight[5][87],
reservoir_weight[5][88],
reservoir_weight[5][89],
reservoir_weight[5][90],
reservoir_weight[5][91],
reservoir_weight[5][92],
reservoir_weight[5][93],
reservoir_weight[5][94],
reservoir_weight[5][95],
reservoir_weight[5][96],
reservoir_weight[5][97],
reservoir_weight[5][98],
reservoir_weight[5][99],
reservoir_weight[5][100],
reservoir_weight[5][101],
reservoir_weight[5][102],
reservoir_weight[5][103],
reservoir_weight[5][104],
reservoir_weight[5][105],
reservoir_weight[5][106],
reservoir_weight[5][107],
reservoir_weight[5][108],
reservoir_weight[5][109],
reservoir_weight[5][110],
reservoir_weight[5][111],
reservoir_weight[5][112],
reservoir_weight[5][113],
reservoir_weight[5][114],
reservoir_weight[5][115],
reservoir_weight[5][116],
reservoir_weight[5][117],
reservoir_weight[5][118],
reservoir_weight[5][119],
reservoir_weight[5][120],
reservoir_weight[5][121],
reservoir_weight[5][122],
reservoir_weight[5][123],
reservoir_weight[5][124],
reservoir_weight[5][125],
reservoir_weight[5][126],
reservoir_weight[5][127],
reservoir_weight[5][128],
reservoir_weight[5][129],
reservoir_weight[5][130],
reservoir_weight[5][131],
reservoir_weight[5][132],
reservoir_weight[5][133],
reservoir_weight[5][134],
reservoir_weight[5][135],
reservoir_weight[5][136],
reservoir_weight[5][137],
reservoir_weight[5][138],
reservoir_weight[5][139],
reservoir_weight[5][140],
reservoir_weight[5][141],
reservoir_weight[5][142],
reservoir_weight[5][143],
reservoir_weight[5][144],
reservoir_weight[5][145],
reservoir_weight[5][146],
reservoir_weight[5][147],
reservoir_weight[5][148],
reservoir_weight[5][149],
reservoir_weight[5][150],
reservoir_weight[5][151],
reservoir_weight[5][152],
reservoir_weight[5][153],
reservoir_weight[5][154],
reservoir_weight[5][155],
reservoir_weight[5][156],
reservoir_weight[5][157],
reservoir_weight[5][158],
reservoir_weight[5][159],
reservoir_weight[5][160],
reservoir_weight[5][161],
reservoir_weight[5][162],
reservoir_weight[5][163],
reservoir_weight[5][164],
reservoir_weight[5][165],
reservoir_weight[5][166],
reservoir_weight[5][167],
reservoir_weight[5][168],
reservoir_weight[5][169],
reservoir_weight[5][170],
reservoir_weight[5][171],
reservoir_weight[5][172],
reservoir_weight[5][173],
reservoir_weight[5][174],
reservoir_weight[5][175],
reservoir_weight[5][176],
reservoir_weight[5][177],
reservoir_weight[5][178],
reservoir_weight[5][179],
reservoir_weight[5][180],
reservoir_weight[5][181],
reservoir_weight[5][182],
reservoir_weight[5][183],
reservoir_weight[5][184],
reservoir_weight[5][185],
reservoir_weight[5][186],
reservoir_weight[5][187],
reservoir_weight[5][188],
reservoir_weight[5][189],
reservoir_weight[5][190],
reservoir_weight[5][191],
reservoir_weight[5][192],
reservoir_weight[5][193],
reservoir_weight[5][194],
reservoir_weight[5][195],
reservoir_weight[5][196],
reservoir_weight[5][197],
reservoir_weight[5][198],
reservoir_weight[5][199]
},
{reservoir_weight[6][0],
reservoir_weight[6][1],
reservoir_weight[6][2],
reservoir_weight[6][3],
reservoir_weight[6][4],
reservoir_weight[6][5],
reservoir_weight[6][6],
reservoir_weight[6][7],
reservoir_weight[6][8],
reservoir_weight[6][9],
reservoir_weight[6][10],
reservoir_weight[6][11],
reservoir_weight[6][12],
reservoir_weight[6][13],
reservoir_weight[6][14],
reservoir_weight[6][15],
reservoir_weight[6][16],
reservoir_weight[6][17],
reservoir_weight[6][18],
reservoir_weight[6][19],
reservoir_weight[6][20],
reservoir_weight[6][21],
reservoir_weight[6][22],
reservoir_weight[6][23],
reservoir_weight[6][24],
reservoir_weight[6][25],
reservoir_weight[6][26],
reservoir_weight[6][27],
reservoir_weight[6][28],
reservoir_weight[6][29],
reservoir_weight[6][30],
reservoir_weight[6][31],
reservoir_weight[6][32],
reservoir_weight[6][33],
reservoir_weight[6][34],
reservoir_weight[6][35],
reservoir_weight[6][36],
reservoir_weight[6][37],
reservoir_weight[6][38],
reservoir_weight[6][39],
reservoir_weight[6][40],
reservoir_weight[6][41],
reservoir_weight[6][42],
reservoir_weight[6][43],
reservoir_weight[6][44],
reservoir_weight[6][45],
reservoir_weight[6][46],
reservoir_weight[6][47],
reservoir_weight[6][48],
reservoir_weight[6][49],
reservoir_weight[6][50],
reservoir_weight[6][51],
reservoir_weight[6][52],
reservoir_weight[6][53],
reservoir_weight[6][54],
reservoir_weight[6][55],
reservoir_weight[6][56],
reservoir_weight[6][57],
reservoir_weight[6][58],
reservoir_weight[6][59],
reservoir_weight[6][60],
reservoir_weight[6][61],
reservoir_weight[6][62],
reservoir_weight[6][63],
reservoir_weight[6][64],
reservoir_weight[6][65],
reservoir_weight[6][66],
reservoir_weight[6][67],
reservoir_weight[6][68],
reservoir_weight[6][69],
reservoir_weight[6][70],
reservoir_weight[6][71],
reservoir_weight[6][72],
reservoir_weight[6][73],
reservoir_weight[6][74],
reservoir_weight[6][75],
reservoir_weight[6][76],
reservoir_weight[6][77],
reservoir_weight[6][78],
reservoir_weight[6][79],
reservoir_weight[6][80],
reservoir_weight[6][81],
reservoir_weight[6][82],
reservoir_weight[6][83],
reservoir_weight[6][84],
reservoir_weight[6][85],
reservoir_weight[6][86],
reservoir_weight[6][87],
reservoir_weight[6][88],
reservoir_weight[6][89],
reservoir_weight[6][90],
reservoir_weight[6][91],
reservoir_weight[6][92],
reservoir_weight[6][93],
reservoir_weight[6][94],
reservoir_weight[6][95],
reservoir_weight[6][96],
reservoir_weight[6][97],
reservoir_weight[6][98],
reservoir_weight[6][99],
reservoir_weight[6][100],
reservoir_weight[6][101],
reservoir_weight[6][102],
reservoir_weight[6][103],
reservoir_weight[6][104],
reservoir_weight[6][105],
reservoir_weight[6][106],
reservoir_weight[6][107],
reservoir_weight[6][108],
reservoir_weight[6][109],
reservoir_weight[6][110],
reservoir_weight[6][111],
reservoir_weight[6][112],
reservoir_weight[6][113],
reservoir_weight[6][114],
reservoir_weight[6][115],
reservoir_weight[6][116],
reservoir_weight[6][117],
reservoir_weight[6][118],
reservoir_weight[6][119],
reservoir_weight[6][120],
reservoir_weight[6][121],
reservoir_weight[6][122],
reservoir_weight[6][123],
reservoir_weight[6][124],
reservoir_weight[6][125],
reservoir_weight[6][126],
reservoir_weight[6][127],
reservoir_weight[6][128],
reservoir_weight[6][129],
reservoir_weight[6][130],
reservoir_weight[6][131],
reservoir_weight[6][132],
reservoir_weight[6][133],
reservoir_weight[6][134],
reservoir_weight[6][135],
reservoir_weight[6][136],
reservoir_weight[6][137],
reservoir_weight[6][138],
reservoir_weight[6][139],
reservoir_weight[6][140],
reservoir_weight[6][141],
reservoir_weight[6][142],
reservoir_weight[6][143],
reservoir_weight[6][144],
reservoir_weight[6][145],
reservoir_weight[6][146],
reservoir_weight[6][147],
reservoir_weight[6][148],
reservoir_weight[6][149],
reservoir_weight[6][150],
reservoir_weight[6][151],
reservoir_weight[6][152],
reservoir_weight[6][153],
reservoir_weight[6][154],
reservoir_weight[6][155],
reservoir_weight[6][156],
reservoir_weight[6][157],
reservoir_weight[6][158],
reservoir_weight[6][159],
reservoir_weight[6][160],
reservoir_weight[6][161],
reservoir_weight[6][162],
reservoir_weight[6][163],
reservoir_weight[6][164],
reservoir_weight[6][165],
reservoir_weight[6][166],
reservoir_weight[6][167],
reservoir_weight[6][168],
reservoir_weight[6][169],
reservoir_weight[6][170],
reservoir_weight[6][171],
reservoir_weight[6][172],
reservoir_weight[6][173],
reservoir_weight[6][174],
reservoir_weight[6][175],
reservoir_weight[6][176],
reservoir_weight[6][177],
reservoir_weight[6][178],
reservoir_weight[6][179],
reservoir_weight[6][180],
reservoir_weight[6][181],
reservoir_weight[6][182],
reservoir_weight[6][183],
reservoir_weight[6][184],
reservoir_weight[6][185],
reservoir_weight[6][186],
reservoir_weight[6][187],
reservoir_weight[6][188],
reservoir_weight[6][189],
reservoir_weight[6][190],
reservoir_weight[6][191],
reservoir_weight[6][192],
reservoir_weight[6][193],
reservoir_weight[6][194],
reservoir_weight[6][195],
reservoir_weight[6][196],
reservoir_weight[6][197],
reservoir_weight[6][198],
reservoir_weight[6][199]
},
{reservoir_weight[7][0],
reservoir_weight[7][1],
reservoir_weight[7][2],
reservoir_weight[7][3],
reservoir_weight[7][4],
reservoir_weight[7][5],
reservoir_weight[7][6],
reservoir_weight[7][7],
reservoir_weight[7][8],
reservoir_weight[7][9],
reservoir_weight[7][10],
reservoir_weight[7][11],
reservoir_weight[7][12],
reservoir_weight[7][13],
reservoir_weight[7][14],
reservoir_weight[7][15],
reservoir_weight[7][16],
reservoir_weight[7][17],
reservoir_weight[7][18],
reservoir_weight[7][19],
reservoir_weight[7][20],
reservoir_weight[7][21],
reservoir_weight[7][22],
reservoir_weight[7][23],
reservoir_weight[7][24],
reservoir_weight[7][25],
reservoir_weight[7][26],
reservoir_weight[7][27],
reservoir_weight[7][28],
reservoir_weight[7][29],
reservoir_weight[7][30],
reservoir_weight[7][31],
reservoir_weight[7][32],
reservoir_weight[7][33],
reservoir_weight[7][34],
reservoir_weight[7][35],
reservoir_weight[7][36],
reservoir_weight[7][37],
reservoir_weight[7][38],
reservoir_weight[7][39],
reservoir_weight[7][40],
reservoir_weight[7][41],
reservoir_weight[7][42],
reservoir_weight[7][43],
reservoir_weight[7][44],
reservoir_weight[7][45],
reservoir_weight[7][46],
reservoir_weight[7][47],
reservoir_weight[7][48],
reservoir_weight[7][49],
reservoir_weight[7][50],
reservoir_weight[7][51],
reservoir_weight[7][52],
reservoir_weight[7][53],
reservoir_weight[7][54],
reservoir_weight[7][55],
reservoir_weight[7][56],
reservoir_weight[7][57],
reservoir_weight[7][58],
reservoir_weight[7][59],
reservoir_weight[7][60],
reservoir_weight[7][61],
reservoir_weight[7][62],
reservoir_weight[7][63],
reservoir_weight[7][64],
reservoir_weight[7][65],
reservoir_weight[7][66],
reservoir_weight[7][67],
reservoir_weight[7][68],
reservoir_weight[7][69],
reservoir_weight[7][70],
reservoir_weight[7][71],
reservoir_weight[7][72],
reservoir_weight[7][73],
reservoir_weight[7][74],
reservoir_weight[7][75],
reservoir_weight[7][76],
reservoir_weight[7][77],
reservoir_weight[7][78],
reservoir_weight[7][79],
reservoir_weight[7][80],
reservoir_weight[7][81],
reservoir_weight[7][82],
reservoir_weight[7][83],
reservoir_weight[7][84],
reservoir_weight[7][85],
reservoir_weight[7][86],
reservoir_weight[7][87],
reservoir_weight[7][88],
reservoir_weight[7][89],
reservoir_weight[7][90],
reservoir_weight[7][91],
reservoir_weight[7][92],
reservoir_weight[7][93],
reservoir_weight[7][94],
reservoir_weight[7][95],
reservoir_weight[7][96],
reservoir_weight[7][97],
reservoir_weight[7][98],
reservoir_weight[7][99],
reservoir_weight[7][100],
reservoir_weight[7][101],
reservoir_weight[7][102],
reservoir_weight[7][103],
reservoir_weight[7][104],
reservoir_weight[7][105],
reservoir_weight[7][106],
reservoir_weight[7][107],
reservoir_weight[7][108],
reservoir_weight[7][109],
reservoir_weight[7][110],
reservoir_weight[7][111],
reservoir_weight[7][112],
reservoir_weight[7][113],
reservoir_weight[7][114],
reservoir_weight[7][115],
reservoir_weight[7][116],
reservoir_weight[7][117],
reservoir_weight[7][118],
reservoir_weight[7][119],
reservoir_weight[7][120],
reservoir_weight[7][121],
reservoir_weight[7][122],
reservoir_weight[7][123],
reservoir_weight[7][124],
reservoir_weight[7][125],
reservoir_weight[7][126],
reservoir_weight[7][127],
reservoir_weight[7][128],
reservoir_weight[7][129],
reservoir_weight[7][130],
reservoir_weight[7][131],
reservoir_weight[7][132],
reservoir_weight[7][133],
reservoir_weight[7][134],
reservoir_weight[7][135],
reservoir_weight[7][136],
reservoir_weight[7][137],
reservoir_weight[7][138],
reservoir_weight[7][139],
reservoir_weight[7][140],
reservoir_weight[7][141],
reservoir_weight[7][142],
reservoir_weight[7][143],
reservoir_weight[7][144],
reservoir_weight[7][145],
reservoir_weight[7][146],
reservoir_weight[7][147],
reservoir_weight[7][148],
reservoir_weight[7][149],
reservoir_weight[7][150],
reservoir_weight[7][151],
reservoir_weight[7][152],
reservoir_weight[7][153],
reservoir_weight[7][154],
reservoir_weight[7][155],
reservoir_weight[7][156],
reservoir_weight[7][157],
reservoir_weight[7][158],
reservoir_weight[7][159],
reservoir_weight[7][160],
reservoir_weight[7][161],
reservoir_weight[7][162],
reservoir_weight[7][163],
reservoir_weight[7][164],
reservoir_weight[7][165],
reservoir_weight[7][166],
reservoir_weight[7][167],
reservoir_weight[7][168],
reservoir_weight[7][169],
reservoir_weight[7][170],
reservoir_weight[7][171],
reservoir_weight[7][172],
reservoir_weight[7][173],
reservoir_weight[7][174],
reservoir_weight[7][175],
reservoir_weight[7][176],
reservoir_weight[7][177],
reservoir_weight[7][178],
reservoir_weight[7][179],
reservoir_weight[7][180],
reservoir_weight[7][181],
reservoir_weight[7][182],
reservoir_weight[7][183],
reservoir_weight[7][184],
reservoir_weight[7][185],
reservoir_weight[7][186],
reservoir_weight[7][187],
reservoir_weight[7][188],
reservoir_weight[7][189],
reservoir_weight[7][190],
reservoir_weight[7][191],
reservoir_weight[7][192],
reservoir_weight[7][193],
reservoir_weight[7][194],
reservoir_weight[7][195],
reservoir_weight[7][196],
reservoir_weight[7][197],
reservoir_weight[7][198],
reservoir_weight[7][199]
},
{reservoir_weight[8][0],
reservoir_weight[8][1],
reservoir_weight[8][2],
reservoir_weight[8][3],
reservoir_weight[8][4],
reservoir_weight[8][5],
reservoir_weight[8][6],
reservoir_weight[8][7],
reservoir_weight[8][8],
reservoir_weight[8][9],
reservoir_weight[8][10],
reservoir_weight[8][11],
reservoir_weight[8][12],
reservoir_weight[8][13],
reservoir_weight[8][14],
reservoir_weight[8][15],
reservoir_weight[8][16],
reservoir_weight[8][17],
reservoir_weight[8][18],
reservoir_weight[8][19],
reservoir_weight[8][20],
reservoir_weight[8][21],
reservoir_weight[8][22],
reservoir_weight[8][23],
reservoir_weight[8][24],
reservoir_weight[8][25],
reservoir_weight[8][26],
reservoir_weight[8][27],
reservoir_weight[8][28],
reservoir_weight[8][29],
reservoir_weight[8][30],
reservoir_weight[8][31],
reservoir_weight[8][32],
reservoir_weight[8][33],
reservoir_weight[8][34],
reservoir_weight[8][35],
reservoir_weight[8][36],
reservoir_weight[8][37],
reservoir_weight[8][38],
reservoir_weight[8][39],
reservoir_weight[8][40],
reservoir_weight[8][41],
reservoir_weight[8][42],
reservoir_weight[8][43],
reservoir_weight[8][44],
reservoir_weight[8][45],
reservoir_weight[8][46],
reservoir_weight[8][47],
reservoir_weight[8][48],
reservoir_weight[8][49],
reservoir_weight[8][50],
reservoir_weight[8][51],
reservoir_weight[8][52],
reservoir_weight[8][53],
reservoir_weight[8][54],
reservoir_weight[8][55],
reservoir_weight[8][56],
reservoir_weight[8][57],
reservoir_weight[8][58],
reservoir_weight[8][59],
reservoir_weight[8][60],
reservoir_weight[8][61],
reservoir_weight[8][62],
reservoir_weight[8][63],
reservoir_weight[8][64],
reservoir_weight[8][65],
reservoir_weight[8][66],
reservoir_weight[8][67],
reservoir_weight[8][68],
reservoir_weight[8][69],
reservoir_weight[8][70],
reservoir_weight[8][71],
reservoir_weight[8][72],
reservoir_weight[8][73],
reservoir_weight[8][74],
reservoir_weight[8][75],
reservoir_weight[8][76],
reservoir_weight[8][77],
reservoir_weight[8][78],
reservoir_weight[8][79],
reservoir_weight[8][80],
reservoir_weight[8][81],
reservoir_weight[8][82],
reservoir_weight[8][83],
reservoir_weight[8][84],
reservoir_weight[8][85],
reservoir_weight[8][86],
reservoir_weight[8][87],
reservoir_weight[8][88],
reservoir_weight[8][89],
reservoir_weight[8][90],
reservoir_weight[8][91],
reservoir_weight[8][92],
reservoir_weight[8][93],
reservoir_weight[8][94],
reservoir_weight[8][95],
reservoir_weight[8][96],
reservoir_weight[8][97],
reservoir_weight[8][98],
reservoir_weight[8][99],
reservoir_weight[8][100],
reservoir_weight[8][101],
reservoir_weight[8][102],
reservoir_weight[8][103],
reservoir_weight[8][104],
reservoir_weight[8][105],
reservoir_weight[8][106],
reservoir_weight[8][107],
reservoir_weight[8][108],
reservoir_weight[8][109],
reservoir_weight[8][110],
reservoir_weight[8][111],
reservoir_weight[8][112],
reservoir_weight[8][113],
reservoir_weight[8][114],
reservoir_weight[8][115],
reservoir_weight[8][116],
reservoir_weight[8][117],
reservoir_weight[8][118],
reservoir_weight[8][119],
reservoir_weight[8][120],
reservoir_weight[8][121],
reservoir_weight[8][122],
reservoir_weight[8][123],
reservoir_weight[8][124],
reservoir_weight[8][125],
reservoir_weight[8][126],
reservoir_weight[8][127],
reservoir_weight[8][128],
reservoir_weight[8][129],
reservoir_weight[8][130],
reservoir_weight[8][131],
reservoir_weight[8][132],
reservoir_weight[8][133],
reservoir_weight[8][134],
reservoir_weight[8][135],
reservoir_weight[8][136],
reservoir_weight[8][137],
reservoir_weight[8][138],
reservoir_weight[8][139],
reservoir_weight[8][140],
reservoir_weight[8][141],
reservoir_weight[8][142],
reservoir_weight[8][143],
reservoir_weight[8][144],
reservoir_weight[8][145],
reservoir_weight[8][146],
reservoir_weight[8][147],
reservoir_weight[8][148],
reservoir_weight[8][149],
reservoir_weight[8][150],
reservoir_weight[8][151],
reservoir_weight[8][152],
reservoir_weight[8][153],
reservoir_weight[8][154],
reservoir_weight[8][155],
reservoir_weight[8][156],
reservoir_weight[8][157],
reservoir_weight[8][158],
reservoir_weight[8][159],
reservoir_weight[8][160],
reservoir_weight[8][161],
reservoir_weight[8][162],
reservoir_weight[8][163],
reservoir_weight[8][164],
reservoir_weight[8][165],
reservoir_weight[8][166],
reservoir_weight[8][167],
reservoir_weight[8][168],
reservoir_weight[8][169],
reservoir_weight[8][170],
reservoir_weight[8][171],
reservoir_weight[8][172],
reservoir_weight[8][173],
reservoir_weight[8][174],
reservoir_weight[8][175],
reservoir_weight[8][176],
reservoir_weight[8][177],
reservoir_weight[8][178],
reservoir_weight[8][179],
reservoir_weight[8][180],
reservoir_weight[8][181],
reservoir_weight[8][182],
reservoir_weight[8][183],
reservoir_weight[8][184],
reservoir_weight[8][185],
reservoir_weight[8][186],
reservoir_weight[8][187],
reservoir_weight[8][188],
reservoir_weight[8][189],
reservoir_weight[8][190],
reservoir_weight[8][191],
reservoir_weight[8][192],
reservoir_weight[8][193],
reservoir_weight[8][194],
reservoir_weight[8][195],
reservoir_weight[8][196],
reservoir_weight[8][197],
reservoir_weight[8][198],
reservoir_weight[8][199]
},
{reservoir_weight[9][0],
reservoir_weight[9][1],
reservoir_weight[9][2],
reservoir_weight[9][3],
reservoir_weight[9][4],
reservoir_weight[9][5],
reservoir_weight[9][6],
reservoir_weight[9][7],
reservoir_weight[9][8],
reservoir_weight[9][9],
reservoir_weight[9][10],
reservoir_weight[9][11],
reservoir_weight[9][12],
reservoir_weight[9][13],
reservoir_weight[9][14],
reservoir_weight[9][15],
reservoir_weight[9][16],
reservoir_weight[9][17],
reservoir_weight[9][18],
reservoir_weight[9][19],
reservoir_weight[9][20],
reservoir_weight[9][21],
reservoir_weight[9][22],
reservoir_weight[9][23],
reservoir_weight[9][24],
reservoir_weight[9][25],
reservoir_weight[9][26],
reservoir_weight[9][27],
reservoir_weight[9][28],
reservoir_weight[9][29],
reservoir_weight[9][30],
reservoir_weight[9][31],
reservoir_weight[9][32],
reservoir_weight[9][33],
reservoir_weight[9][34],
reservoir_weight[9][35],
reservoir_weight[9][36],
reservoir_weight[9][37],
reservoir_weight[9][38],
reservoir_weight[9][39],
reservoir_weight[9][40],
reservoir_weight[9][41],
reservoir_weight[9][42],
reservoir_weight[9][43],
reservoir_weight[9][44],
reservoir_weight[9][45],
reservoir_weight[9][46],
reservoir_weight[9][47],
reservoir_weight[9][48],
reservoir_weight[9][49],
reservoir_weight[9][50],
reservoir_weight[9][51],
reservoir_weight[9][52],
reservoir_weight[9][53],
reservoir_weight[9][54],
reservoir_weight[9][55],
reservoir_weight[9][56],
reservoir_weight[9][57],
reservoir_weight[9][58],
reservoir_weight[9][59],
reservoir_weight[9][60],
reservoir_weight[9][61],
reservoir_weight[9][62],
reservoir_weight[9][63],
reservoir_weight[9][64],
reservoir_weight[9][65],
reservoir_weight[9][66],
reservoir_weight[9][67],
reservoir_weight[9][68],
reservoir_weight[9][69],
reservoir_weight[9][70],
reservoir_weight[9][71],
reservoir_weight[9][72],
reservoir_weight[9][73],
reservoir_weight[9][74],
reservoir_weight[9][75],
reservoir_weight[9][76],
reservoir_weight[9][77],
reservoir_weight[9][78],
reservoir_weight[9][79],
reservoir_weight[9][80],
reservoir_weight[9][81],
reservoir_weight[9][82],
reservoir_weight[9][83],
reservoir_weight[9][84],
reservoir_weight[9][85],
reservoir_weight[9][86],
reservoir_weight[9][87],
reservoir_weight[9][88],
reservoir_weight[9][89],
reservoir_weight[9][90],
reservoir_weight[9][91],
reservoir_weight[9][92],
reservoir_weight[9][93],
reservoir_weight[9][94],
reservoir_weight[9][95],
reservoir_weight[9][96],
reservoir_weight[9][97],
reservoir_weight[9][98],
reservoir_weight[9][99],
reservoir_weight[9][100],
reservoir_weight[9][101],
reservoir_weight[9][102],
reservoir_weight[9][103],
reservoir_weight[9][104],
reservoir_weight[9][105],
reservoir_weight[9][106],
reservoir_weight[9][107],
reservoir_weight[9][108],
reservoir_weight[9][109],
reservoir_weight[9][110],
reservoir_weight[9][111],
reservoir_weight[9][112],
reservoir_weight[9][113],
reservoir_weight[9][114],
reservoir_weight[9][115],
reservoir_weight[9][116],
reservoir_weight[9][117],
reservoir_weight[9][118],
reservoir_weight[9][119],
reservoir_weight[9][120],
reservoir_weight[9][121],
reservoir_weight[9][122],
reservoir_weight[9][123],
reservoir_weight[9][124],
reservoir_weight[9][125],
reservoir_weight[9][126],
reservoir_weight[9][127],
reservoir_weight[9][128],
reservoir_weight[9][129],
reservoir_weight[9][130],
reservoir_weight[9][131],
reservoir_weight[9][132],
reservoir_weight[9][133],
reservoir_weight[9][134],
reservoir_weight[9][135],
reservoir_weight[9][136],
reservoir_weight[9][137],
reservoir_weight[9][138],
reservoir_weight[9][139],
reservoir_weight[9][140],
reservoir_weight[9][141],
reservoir_weight[9][142],
reservoir_weight[9][143],
reservoir_weight[9][144],
reservoir_weight[9][145],
reservoir_weight[9][146],
reservoir_weight[9][147],
reservoir_weight[9][148],
reservoir_weight[9][149],
reservoir_weight[9][150],
reservoir_weight[9][151],
reservoir_weight[9][152],
reservoir_weight[9][153],
reservoir_weight[9][154],
reservoir_weight[9][155],
reservoir_weight[9][156],
reservoir_weight[9][157],
reservoir_weight[9][158],
reservoir_weight[9][159],
reservoir_weight[9][160],
reservoir_weight[9][161],
reservoir_weight[9][162],
reservoir_weight[9][163],
reservoir_weight[9][164],
reservoir_weight[9][165],
reservoir_weight[9][166],
reservoir_weight[9][167],
reservoir_weight[9][168],
reservoir_weight[9][169],
reservoir_weight[9][170],
reservoir_weight[9][171],
reservoir_weight[9][172],
reservoir_weight[9][173],
reservoir_weight[9][174],
reservoir_weight[9][175],
reservoir_weight[9][176],
reservoir_weight[9][177],
reservoir_weight[9][178],
reservoir_weight[9][179],
reservoir_weight[9][180],
reservoir_weight[9][181],
reservoir_weight[9][182],
reservoir_weight[9][183],
reservoir_weight[9][184],
reservoir_weight[9][185],
reservoir_weight[9][186],
reservoir_weight[9][187],
reservoir_weight[9][188],
reservoir_weight[9][189],
reservoir_weight[9][190],
reservoir_weight[9][191],
reservoir_weight[9][192],
reservoir_weight[9][193],
reservoir_weight[9][194],
reservoir_weight[9][195],
reservoir_weight[9][196],
reservoir_weight[9][197],
reservoir_weight[9][198],
reservoir_weight[9][199]
},
{reservoir_weight[10][0],
reservoir_weight[10][1],
reservoir_weight[10][2],
reservoir_weight[10][3],
reservoir_weight[10][4],
reservoir_weight[10][5],
reservoir_weight[10][6],
reservoir_weight[10][7],
reservoir_weight[10][8],
reservoir_weight[10][9],
reservoir_weight[10][10],
reservoir_weight[10][11],
reservoir_weight[10][12],
reservoir_weight[10][13],
reservoir_weight[10][14],
reservoir_weight[10][15],
reservoir_weight[10][16],
reservoir_weight[10][17],
reservoir_weight[10][18],
reservoir_weight[10][19],
reservoir_weight[10][20],
reservoir_weight[10][21],
reservoir_weight[10][22],
reservoir_weight[10][23],
reservoir_weight[10][24],
reservoir_weight[10][25],
reservoir_weight[10][26],
reservoir_weight[10][27],
reservoir_weight[10][28],
reservoir_weight[10][29],
reservoir_weight[10][30],
reservoir_weight[10][31],
reservoir_weight[10][32],
reservoir_weight[10][33],
reservoir_weight[10][34],
reservoir_weight[10][35],
reservoir_weight[10][36],
reservoir_weight[10][37],
reservoir_weight[10][38],
reservoir_weight[10][39],
reservoir_weight[10][40],
reservoir_weight[10][41],
reservoir_weight[10][42],
reservoir_weight[10][43],
reservoir_weight[10][44],
reservoir_weight[10][45],
reservoir_weight[10][46],
reservoir_weight[10][47],
reservoir_weight[10][48],
reservoir_weight[10][49],
reservoir_weight[10][50],
reservoir_weight[10][51],
reservoir_weight[10][52],
reservoir_weight[10][53],
reservoir_weight[10][54],
reservoir_weight[10][55],
reservoir_weight[10][56],
reservoir_weight[10][57],
reservoir_weight[10][58],
reservoir_weight[10][59],
reservoir_weight[10][60],
reservoir_weight[10][61],
reservoir_weight[10][62],
reservoir_weight[10][63],
reservoir_weight[10][64],
reservoir_weight[10][65],
reservoir_weight[10][66],
reservoir_weight[10][67],
reservoir_weight[10][68],
reservoir_weight[10][69],
reservoir_weight[10][70],
reservoir_weight[10][71],
reservoir_weight[10][72],
reservoir_weight[10][73],
reservoir_weight[10][74],
reservoir_weight[10][75],
reservoir_weight[10][76],
reservoir_weight[10][77],
reservoir_weight[10][78],
reservoir_weight[10][79],
reservoir_weight[10][80],
reservoir_weight[10][81],
reservoir_weight[10][82],
reservoir_weight[10][83],
reservoir_weight[10][84],
reservoir_weight[10][85],
reservoir_weight[10][86],
reservoir_weight[10][87],
reservoir_weight[10][88],
reservoir_weight[10][89],
reservoir_weight[10][90],
reservoir_weight[10][91],
reservoir_weight[10][92],
reservoir_weight[10][93],
reservoir_weight[10][94],
reservoir_weight[10][95],
reservoir_weight[10][96],
reservoir_weight[10][97],
reservoir_weight[10][98],
reservoir_weight[10][99],
reservoir_weight[10][100],
reservoir_weight[10][101],
reservoir_weight[10][102],
reservoir_weight[10][103],
reservoir_weight[10][104],
reservoir_weight[10][105],
reservoir_weight[10][106],
reservoir_weight[10][107],
reservoir_weight[10][108],
reservoir_weight[10][109],
reservoir_weight[10][110],
reservoir_weight[10][111],
reservoir_weight[10][112],
reservoir_weight[10][113],
reservoir_weight[10][114],
reservoir_weight[10][115],
reservoir_weight[10][116],
reservoir_weight[10][117],
reservoir_weight[10][118],
reservoir_weight[10][119],
reservoir_weight[10][120],
reservoir_weight[10][121],
reservoir_weight[10][122],
reservoir_weight[10][123],
reservoir_weight[10][124],
reservoir_weight[10][125],
reservoir_weight[10][126],
reservoir_weight[10][127],
reservoir_weight[10][128],
reservoir_weight[10][129],
reservoir_weight[10][130],
reservoir_weight[10][131],
reservoir_weight[10][132],
reservoir_weight[10][133],
reservoir_weight[10][134],
reservoir_weight[10][135],
reservoir_weight[10][136],
reservoir_weight[10][137],
reservoir_weight[10][138],
reservoir_weight[10][139],
reservoir_weight[10][140],
reservoir_weight[10][141],
reservoir_weight[10][142],
reservoir_weight[10][143],
reservoir_weight[10][144],
reservoir_weight[10][145],
reservoir_weight[10][146],
reservoir_weight[10][147],
reservoir_weight[10][148],
reservoir_weight[10][149],
reservoir_weight[10][150],
reservoir_weight[10][151],
reservoir_weight[10][152],
reservoir_weight[10][153],
reservoir_weight[10][154],
reservoir_weight[10][155],
reservoir_weight[10][156],
reservoir_weight[10][157],
reservoir_weight[10][158],
reservoir_weight[10][159],
reservoir_weight[10][160],
reservoir_weight[10][161],
reservoir_weight[10][162],
reservoir_weight[10][163],
reservoir_weight[10][164],
reservoir_weight[10][165],
reservoir_weight[10][166],
reservoir_weight[10][167],
reservoir_weight[10][168],
reservoir_weight[10][169],
reservoir_weight[10][170],
reservoir_weight[10][171],
reservoir_weight[10][172],
reservoir_weight[10][173],
reservoir_weight[10][174],
reservoir_weight[10][175],
reservoir_weight[10][176],
reservoir_weight[10][177],
reservoir_weight[10][178],
reservoir_weight[10][179],
reservoir_weight[10][180],
reservoir_weight[10][181],
reservoir_weight[10][182],
reservoir_weight[10][183],
reservoir_weight[10][184],
reservoir_weight[10][185],
reservoir_weight[10][186],
reservoir_weight[10][187],
reservoir_weight[10][188],
reservoir_weight[10][189],
reservoir_weight[10][190],
reservoir_weight[10][191],
reservoir_weight[10][192],
reservoir_weight[10][193],
reservoir_weight[10][194],
reservoir_weight[10][195],
reservoir_weight[10][196],
reservoir_weight[10][197],
reservoir_weight[10][198],
reservoir_weight[10][199]
},
{reservoir_weight[11][0],
reservoir_weight[11][1],
reservoir_weight[11][2],
reservoir_weight[11][3],
reservoir_weight[11][4],
reservoir_weight[11][5],
reservoir_weight[11][6],
reservoir_weight[11][7],
reservoir_weight[11][8],
reservoir_weight[11][9],
reservoir_weight[11][10],
reservoir_weight[11][11],
reservoir_weight[11][12],
reservoir_weight[11][13],
reservoir_weight[11][14],
reservoir_weight[11][15],
reservoir_weight[11][16],
reservoir_weight[11][17],
reservoir_weight[11][18],
reservoir_weight[11][19],
reservoir_weight[11][20],
reservoir_weight[11][21],
reservoir_weight[11][22],
reservoir_weight[11][23],
reservoir_weight[11][24],
reservoir_weight[11][25],
reservoir_weight[11][26],
reservoir_weight[11][27],
reservoir_weight[11][28],
reservoir_weight[11][29],
reservoir_weight[11][30],
reservoir_weight[11][31],
reservoir_weight[11][32],
reservoir_weight[11][33],
reservoir_weight[11][34],
reservoir_weight[11][35],
reservoir_weight[11][36],
reservoir_weight[11][37],
reservoir_weight[11][38],
reservoir_weight[11][39],
reservoir_weight[11][40],
reservoir_weight[11][41],
reservoir_weight[11][42],
reservoir_weight[11][43],
reservoir_weight[11][44],
reservoir_weight[11][45],
reservoir_weight[11][46],
reservoir_weight[11][47],
reservoir_weight[11][48],
reservoir_weight[11][49],
reservoir_weight[11][50],
reservoir_weight[11][51],
reservoir_weight[11][52],
reservoir_weight[11][53],
reservoir_weight[11][54],
reservoir_weight[11][55],
reservoir_weight[11][56],
reservoir_weight[11][57],
reservoir_weight[11][58],
reservoir_weight[11][59],
reservoir_weight[11][60],
reservoir_weight[11][61],
reservoir_weight[11][62],
reservoir_weight[11][63],
reservoir_weight[11][64],
reservoir_weight[11][65],
reservoir_weight[11][66],
reservoir_weight[11][67],
reservoir_weight[11][68],
reservoir_weight[11][69],
reservoir_weight[11][70],
reservoir_weight[11][71],
reservoir_weight[11][72],
reservoir_weight[11][73],
reservoir_weight[11][74],
reservoir_weight[11][75],
reservoir_weight[11][76],
reservoir_weight[11][77],
reservoir_weight[11][78],
reservoir_weight[11][79],
reservoir_weight[11][80],
reservoir_weight[11][81],
reservoir_weight[11][82],
reservoir_weight[11][83],
reservoir_weight[11][84],
reservoir_weight[11][85],
reservoir_weight[11][86],
reservoir_weight[11][87],
reservoir_weight[11][88],
reservoir_weight[11][89],
reservoir_weight[11][90],
reservoir_weight[11][91],
reservoir_weight[11][92],
reservoir_weight[11][93],
reservoir_weight[11][94],
reservoir_weight[11][95],
reservoir_weight[11][96],
reservoir_weight[11][97],
reservoir_weight[11][98],
reservoir_weight[11][99],
reservoir_weight[11][100],
reservoir_weight[11][101],
reservoir_weight[11][102],
reservoir_weight[11][103],
reservoir_weight[11][104],
reservoir_weight[11][105],
reservoir_weight[11][106],
reservoir_weight[11][107],
reservoir_weight[11][108],
reservoir_weight[11][109],
reservoir_weight[11][110],
reservoir_weight[11][111],
reservoir_weight[11][112],
reservoir_weight[11][113],
reservoir_weight[11][114],
reservoir_weight[11][115],
reservoir_weight[11][116],
reservoir_weight[11][117],
reservoir_weight[11][118],
reservoir_weight[11][119],
reservoir_weight[11][120],
reservoir_weight[11][121],
reservoir_weight[11][122],
reservoir_weight[11][123],
reservoir_weight[11][124],
reservoir_weight[11][125],
reservoir_weight[11][126],
reservoir_weight[11][127],
reservoir_weight[11][128],
reservoir_weight[11][129],
reservoir_weight[11][130],
reservoir_weight[11][131],
reservoir_weight[11][132],
reservoir_weight[11][133],
reservoir_weight[11][134],
reservoir_weight[11][135],
reservoir_weight[11][136],
reservoir_weight[11][137],
reservoir_weight[11][138],
reservoir_weight[11][139],
reservoir_weight[11][140],
reservoir_weight[11][141],
reservoir_weight[11][142],
reservoir_weight[11][143],
reservoir_weight[11][144],
reservoir_weight[11][145],
reservoir_weight[11][146],
reservoir_weight[11][147],
reservoir_weight[11][148],
reservoir_weight[11][149],
reservoir_weight[11][150],
reservoir_weight[11][151],
reservoir_weight[11][152],
reservoir_weight[11][153],
reservoir_weight[11][154],
reservoir_weight[11][155],
reservoir_weight[11][156],
reservoir_weight[11][157],
reservoir_weight[11][158],
reservoir_weight[11][159],
reservoir_weight[11][160],
reservoir_weight[11][161],
reservoir_weight[11][162],
reservoir_weight[11][163],
reservoir_weight[11][164],
reservoir_weight[11][165],
reservoir_weight[11][166],
reservoir_weight[11][167],
reservoir_weight[11][168],
reservoir_weight[11][169],
reservoir_weight[11][170],
reservoir_weight[11][171],
reservoir_weight[11][172],
reservoir_weight[11][173],
reservoir_weight[11][174],
reservoir_weight[11][175],
reservoir_weight[11][176],
reservoir_weight[11][177],
reservoir_weight[11][178],
reservoir_weight[11][179],
reservoir_weight[11][180],
reservoir_weight[11][181],
reservoir_weight[11][182],
reservoir_weight[11][183],
reservoir_weight[11][184],
reservoir_weight[11][185],
reservoir_weight[11][186],
reservoir_weight[11][187],
reservoir_weight[11][188],
reservoir_weight[11][189],
reservoir_weight[11][190],
reservoir_weight[11][191],
reservoir_weight[11][192],
reservoir_weight[11][193],
reservoir_weight[11][194],
reservoir_weight[11][195],
reservoir_weight[11][196],
reservoir_weight[11][197],
reservoir_weight[11][198],
reservoir_weight[11][199]
},
{reservoir_weight[12][0],
reservoir_weight[12][1],
reservoir_weight[12][2],
reservoir_weight[12][3],
reservoir_weight[12][4],
reservoir_weight[12][5],
reservoir_weight[12][6],
reservoir_weight[12][7],
reservoir_weight[12][8],
reservoir_weight[12][9],
reservoir_weight[12][10],
reservoir_weight[12][11],
reservoir_weight[12][12],
reservoir_weight[12][13],
reservoir_weight[12][14],
reservoir_weight[12][15],
reservoir_weight[12][16],
reservoir_weight[12][17],
reservoir_weight[12][18],
reservoir_weight[12][19],
reservoir_weight[12][20],
reservoir_weight[12][21],
reservoir_weight[12][22],
reservoir_weight[12][23],
reservoir_weight[12][24],
reservoir_weight[12][25],
reservoir_weight[12][26],
reservoir_weight[12][27],
reservoir_weight[12][28],
reservoir_weight[12][29],
reservoir_weight[12][30],
reservoir_weight[12][31],
reservoir_weight[12][32],
reservoir_weight[12][33],
reservoir_weight[12][34],
reservoir_weight[12][35],
reservoir_weight[12][36],
reservoir_weight[12][37],
reservoir_weight[12][38],
reservoir_weight[12][39],
reservoir_weight[12][40],
reservoir_weight[12][41],
reservoir_weight[12][42],
reservoir_weight[12][43],
reservoir_weight[12][44],
reservoir_weight[12][45],
reservoir_weight[12][46],
reservoir_weight[12][47],
reservoir_weight[12][48],
reservoir_weight[12][49],
reservoir_weight[12][50],
reservoir_weight[12][51],
reservoir_weight[12][52],
reservoir_weight[12][53],
reservoir_weight[12][54],
reservoir_weight[12][55],
reservoir_weight[12][56],
reservoir_weight[12][57],
reservoir_weight[12][58],
reservoir_weight[12][59],
reservoir_weight[12][60],
reservoir_weight[12][61],
reservoir_weight[12][62],
reservoir_weight[12][63],
reservoir_weight[12][64],
reservoir_weight[12][65],
reservoir_weight[12][66],
reservoir_weight[12][67],
reservoir_weight[12][68],
reservoir_weight[12][69],
reservoir_weight[12][70],
reservoir_weight[12][71],
reservoir_weight[12][72],
reservoir_weight[12][73],
reservoir_weight[12][74],
reservoir_weight[12][75],
reservoir_weight[12][76],
reservoir_weight[12][77],
reservoir_weight[12][78],
reservoir_weight[12][79],
reservoir_weight[12][80],
reservoir_weight[12][81],
reservoir_weight[12][82],
reservoir_weight[12][83],
reservoir_weight[12][84],
reservoir_weight[12][85],
reservoir_weight[12][86],
reservoir_weight[12][87],
reservoir_weight[12][88],
reservoir_weight[12][89],
reservoir_weight[12][90],
reservoir_weight[12][91],
reservoir_weight[12][92],
reservoir_weight[12][93],
reservoir_weight[12][94],
reservoir_weight[12][95],
reservoir_weight[12][96],
reservoir_weight[12][97],
reservoir_weight[12][98],
reservoir_weight[12][99],
reservoir_weight[12][100],
reservoir_weight[12][101],
reservoir_weight[12][102],
reservoir_weight[12][103],
reservoir_weight[12][104],
reservoir_weight[12][105],
reservoir_weight[12][106],
reservoir_weight[12][107],
reservoir_weight[12][108],
reservoir_weight[12][109],
reservoir_weight[12][110],
reservoir_weight[12][111],
reservoir_weight[12][112],
reservoir_weight[12][113],
reservoir_weight[12][114],
reservoir_weight[12][115],
reservoir_weight[12][116],
reservoir_weight[12][117],
reservoir_weight[12][118],
reservoir_weight[12][119],
reservoir_weight[12][120],
reservoir_weight[12][121],
reservoir_weight[12][122],
reservoir_weight[12][123],
reservoir_weight[12][124],
reservoir_weight[12][125],
reservoir_weight[12][126],
reservoir_weight[12][127],
reservoir_weight[12][128],
reservoir_weight[12][129],
reservoir_weight[12][130],
reservoir_weight[12][131],
reservoir_weight[12][132],
reservoir_weight[12][133],
reservoir_weight[12][134],
reservoir_weight[12][135],
reservoir_weight[12][136],
reservoir_weight[12][137],
reservoir_weight[12][138],
reservoir_weight[12][139],
reservoir_weight[12][140],
reservoir_weight[12][141],
reservoir_weight[12][142],
reservoir_weight[12][143],
reservoir_weight[12][144],
reservoir_weight[12][145],
reservoir_weight[12][146],
reservoir_weight[12][147],
reservoir_weight[12][148],
reservoir_weight[12][149],
reservoir_weight[12][150],
reservoir_weight[12][151],
reservoir_weight[12][152],
reservoir_weight[12][153],
reservoir_weight[12][154],
reservoir_weight[12][155],
reservoir_weight[12][156],
reservoir_weight[12][157],
reservoir_weight[12][158],
reservoir_weight[12][159],
reservoir_weight[12][160],
reservoir_weight[12][161],
reservoir_weight[12][162],
reservoir_weight[12][163],
reservoir_weight[12][164],
reservoir_weight[12][165],
reservoir_weight[12][166],
reservoir_weight[12][167],
reservoir_weight[12][168],
reservoir_weight[12][169],
reservoir_weight[12][170],
reservoir_weight[12][171],
reservoir_weight[12][172],
reservoir_weight[12][173],
reservoir_weight[12][174],
reservoir_weight[12][175],
reservoir_weight[12][176],
reservoir_weight[12][177],
reservoir_weight[12][178],
reservoir_weight[12][179],
reservoir_weight[12][180],
reservoir_weight[12][181],
reservoir_weight[12][182],
reservoir_weight[12][183],
reservoir_weight[12][184],
reservoir_weight[12][185],
reservoir_weight[12][186],
reservoir_weight[12][187],
reservoir_weight[12][188],
reservoir_weight[12][189],
reservoir_weight[12][190],
reservoir_weight[12][191],
reservoir_weight[12][192],
reservoir_weight[12][193],
reservoir_weight[12][194],
reservoir_weight[12][195],
reservoir_weight[12][196],
reservoir_weight[12][197],
reservoir_weight[12][198],
reservoir_weight[12][199]
},
{reservoir_weight[13][0],
reservoir_weight[13][1],
reservoir_weight[13][2],
reservoir_weight[13][3],
reservoir_weight[13][4],
reservoir_weight[13][5],
reservoir_weight[13][6],
reservoir_weight[13][7],
reservoir_weight[13][8],
reservoir_weight[13][9],
reservoir_weight[13][10],
reservoir_weight[13][11],
reservoir_weight[13][12],
reservoir_weight[13][13],
reservoir_weight[13][14],
reservoir_weight[13][15],
reservoir_weight[13][16],
reservoir_weight[13][17],
reservoir_weight[13][18],
reservoir_weight[13][19],
reservoir_weight[13][20],
reservoir_weight[13][21],
reservoir_weight[13][22],
reservoir_weight[13][23],
reservoir_weight[13][24],
reservoir_weight[13][25],
reservoir_weight[13][26],
reservoir_weight[13][27],
reservoir_weight[13][28],
reservoir_weight[13][29],
reservoir_weight[13][30],
reservoir_weight[13][31],
reservoir_weight[13][32],
reservoir_weight[13][33],
reservoir_weight[13][34],
reservoir_weight[13][35],
reservoir_weight[13][36],
reservoir_weight[13][37],
reservoir_weight[13][38],
reservoir_weight[13][39],
reservoir_weight[13][40],
reservoir_weight[13][41],
reservoir_weight[13][42],
reservoir_weight[13][43],
reservoir_weight[13][44],
reservoir_weight[13][45],
reservoir_weight[13][46],
reservoir_weight[13][47],
reservoir_weight[13][48],
reservoir_weight[13][49],
reservoir_weight[13][50],
reservoir_weight[13][51],
reservoir_weight[13][52],
reservoir_weight[13][53],
reservoir_weight[13][54],
reservoir_weight[13][55],
reservoir_weight[13][56],
reservoir_weight[13][57],
reservoir_weight[13][58],
reservoir_weight[13][59],
reservoir_weight[13][60],
reservoir_weight[13][61],
reservoir_weight[13][62],
reservoir_weight[13][63],
reservoir_weight[13][64],
reservoir_weight[13][65],
reservoir_weight[13][66],
reservoir_weight[13][67],
reservoir_weight[13][68],
reservoir_weight[13][69],
reservoir_weight[13][70],
reservoir_weight[13][71],
reservoir_weight[13][72],
reservoir_weight[13][73],
reservoir_weight[13][74],
reservoir_weight[13][75],
reservoir_weight[13][76],
reservoir_weight[13][77],
reservoir_weight[13][78],
reservoir_weight[13][79],
reservoir_weight[13][80],
reservoir_weight[13][81],
reservoir_weight[13][82],
reservoir_weight[13][83],
reservoir_weight[13][84],
reservoir_weight[13][85],
reservoir_weight[13][86],
reservoir_weight[13][87],
reservoir_weight[13][88],
reservoir_weight[13][89],
reservoir_weight[13][90],
reservoir_weight[13][91],
reservoir_weight[13][92],
reservoir_weight[13][93],
reservoir_weight[13][94],
reservoir_weight[13][95],
reservoir_weight[13][96],
reservoir_weight[13][97],
reservoir_weight[13][98],
reservoir_weight[13][99],
reservoir_weight[13][100],
reservoir_weight[13][101],
reservoir_weight[13][102],
reservoir_weight[13][103],
reservoir_weight[13][104],
reservoir_weight[13][105],
reservoir_weight[13][106],
reservoir_weight[13][107],
reservoir_weight[13][108],
reservoir_weight[13][109],
reservoir_weight[13][110],
reservoir_weight[13][111],
reservoir_weight[13][112],
reservoir_weight[13][113],
reservoir_weight[13][114],
reservoir_weight[13][115],
reservoir_weight[13][116],
reservoir_weight[13][117],
reservoir_weight[13][118],
reservoir_weight[13][119],
reservoir_weight[13][120],
reservoir_weight[13][121],
reservoir_weight[13][122],
reservoir_weight[13][123],
reservoir_weight[13][124],
reservoir_weight[13][125],
reservoir_weight[13][126],
reservoir_weight[13][127],
reservoir_weight[13][128],
reservoir_weight[13][129],
reservoir_weight[13][130],
reservoir_weight[13][131],
reservoir_weight[13][132],
reservoir_weight[13][133],
reservoir_weight[13][134],
reservoir_weight[13][135],
reservoir_weight[13][136],
reservoir_weight[13][137],
reservoir_weight[13][138],
reservoir_weight[13][139],
reservoir_weight[13][140],
reservoir_weight[13][141],
reservoir_weight[13][142],
reservoir_weight[13][143],
reservoir_weight[13][144],
reservoir_weight[13][145],
reservoir_weight[13][146],
reservoir_weight[13][147],
reservoir_weight[13][148],
reservoir_weight[13][149],
reservoir_weight[13][150],
reservoir_weight[13][151],
reservoir_weight[13][152],
reservoir_weight[13][153],
reservoir_weight[13][154],
reservoir_weight[13][155],
reservoir_weight[13][156],
reservoir_weight[13][157],
reservoir_weight[13][158],
reservoir_weight[13][159],
reservoir_weight[13][160],
reservoir_weight[13][161],
reservoir_weight[13][162],
reservoir_weight[13][163],
reservoir_weight[13][164],
reservoir_weight[13][165],
reservoir_weight[13][166],
reservoir_weight[13][167],
reservoir_weight[13][168],
reservoir_weight[13][169],
reservoir_weight[13][170],
reservoir_weight[13][171],
reservoir_weight[13][172],
reservoir_weight[13][173],
reservoir_weight[13][174],
reservoir_weight[13][175],
reservoir_weight[13][176],
reservoir_weight[13][177],
reservoir_weight[13][178],
reservoir_weight[13][179],
reservoir_weight[13][180],
reservoir_weight[13][181],
reservoir_weight[13][182],
reservoir_weight[13][183],
reservoir_weight[13][184],
reservoir_weight[13][185],
reservoir_weight[13][186],
reservoir_weight[13][187],
reservoir_weight[13][188],
reservoir_weight[13][189],
reservoir_weight[13][190],
reservoir_weight[13][191],
reservoir_weight[13][192],
reservoir_weight[13][193],
reservoir_weight[13][194],
reservoir_weight[13][195],
reservoir_weight[13][196],
reservoir_weight[13][197],
reservoir_weight[13][198],
reservoir_weight[13][199]
},
{reservoir_weight[14][0],
reservoir_weight[14][1],
reservoir_weight[14][2],
reservoir_weight[14][3],
reservoir_weight[14][4],
reservoir_weight[14][5],
reservoir_weight[14][6],
reservoir_weight[14][7],
reservoir_weight[14][8],
reservoir_weight[14][9],
reservoir_weight[14][10],
reservoir_weight[14][11],
reservoir_weight[14][12],
reservoir_weight[14][13],
reservoir_weight[14][14],
reservoir_weight[14][15],
reservoir_weight[14][16],
reservoir_weight[14][17],
reservoir_weight[14][18],
reservoir_weight[14][19],
reservoir_weight[14][20],
reservoir_weight[14][21],
reservoir_weight[14][22],
reservoir_weight[14][23],
reservoir_weight[14][24],
reservoir_weight[14][25],
reservoir_weight[14][26],
reservoir_weight[14][27],
reservoir_weight[14][28],
reservoir_weight[14][29],
reservoir_weight[14][30],
reservoir_weight[14][31],
reservoir_weight[14][32],
reservoir_weight[14][33],
reservoir_weight[14][34],
reservoir_weight[14][35],
reservoir_weight[14][36],
reservoir_weight[14][37],
reservoir_weight[14][38],
reservoir_weight[14][39],
reservoir_weight[14][40],
reservoir_weight[14][41],
reservoir_weight[14][42],
reservoir_weight[14][43],
reservoir_weight[14][44],
reservoir_weight[14][45],
reservoir_weight[14][46],
reservoir_weight[14][47],
reservoir_weight[14][48],
reservoir_weight[14][49],
reservoir_weight[14][50],
reservoir_weight[14][51],
reservoir_weight[14][52],
reservoir_weight[14][53],
reservoir_weight[14][54],
reservoir_weight[14][55],
reservoir_weight[14][56],
reservoir_weight[14][57],
reservoir_weight[14][58],
reservoir_weight[14][59],
reservoir_weight[14][60],
reservoir_weight[14][61],
reservoir_weight[14][62],
reservoir_weight[14][63],
reservoir_weight[14][64],
reservoir_weight[14][65],
reservoir_weight[14][66],
reservoir_weight[14][67],
reservoir_weight[14][68],
reservoir_weight[14][69],
reservoir_weight[14][70],
reservoir_weight[14][71],
reservoir_weight[14][72],
reservoir_weight[14][73],
reservoir_weight[14][74],
reservoir_weight[14][75],
reservoir_weight[14][76],
reservoir_weight[14][77],
reservoir_weight[14][78],
reservoir_weight[14][79],
reservoir_weight[14][80],
reservoir_weight[14][81],
reservoir_weight[14][82],
reservoir_weight[14][83],
reservoir_weight[14][84],
reservoir_weight[14][85],
reservoir_weight[14][86],
reservoir_weight[14][87],
reservoir_weight[14][88],
reservoir_weight[14][89],
reservoir_weight[14][90],
reservoir_weight[14][91],
reservoir_weight[14][92],
reservoir_weight[14][93],
reservoir_weight[14][94],
reservoir_weight[14][95],
reservoir_weight[14][96],
reservoir_weight[14][97],
reservoir_weight[14][98],
reservoir_weight[14][99],
reservoir_weight[14][100],
reservoir_weight[14][101],
reservoir_weight[14][102],
reservoir_weight[14][103],
reservoir_weight[14][104],
reservoir_weight[14][105],
reservoir_weight[14][106],
reservoir_weight[14][107],
reservoir_weight[14][108],
reservoir_weight[14][109],
reservoir_weight[14][110],
reservoir_weight[14][111],
reservoir_weight[14][112],
reservoir_weight[14][113],
reservoir_weight[14][114],
reservoir_weight[14][115],
reservoir_weight[14][116],
reservoir_weight[14][117],
reservoir_weight[14][118],
reservoir_weight[14][119],
reservoir_weight[14][120],
reservoir_weight[14][121],
reservoir_weight[14][122],
reservoir_weight[14][123],
reservoir_weight[14][124],
reservoir_weight[14][125],
reservoir_weight[14][126],
reservoir_weight[14][127],
reservoir_weight[14][128],
reservoir_weight[14][129],
reservoir_weight[14][130],
reservoir_weight[14][131],
reservoir_weight[14][132],
reservoir_weight[14][133],
reservoir_weight[14][134],
reservoir_weight[14][135],
reservoir_weight[14][136],
reservoir_weight[14][137],
reservoir_weight[14][138],
reservoir_weight[14][139],
reservoir_weight[14][140],
reservoir_weight[14][141],
reservoir_weight[14][142],
reservoir_weight[14][143],
reservoir_weight[14][144],
reservoir_weight[14][145],
reservoir_weight[14][146],
reservoir_weight[14][147],
reservoir_weight[14][148],
reservoir_weight[14][149],
reservoir_weight[14][150],
reservoir_weight[14][151],
reservoir_weight[14][152],
reservoir_weight[14][153],
reservoir_weight[14][154],
reservoir_weight[14][155],
reservoir_weight[14][156],
reservoir_weight[14][157],
reservoir_weight[14][158],
reservoir_weight[14][159],
reservoir_weight[14][160],
reservoir_weight[14][161],
reservoir_weight[14][162],
reservoir_weight[14][163],
reservoir_weight[14][164],
reservoir_weight[14][165],
reservoir_weight[14][166],
reservoir_weight[14][167],
reservoir_weight[14][168],
reservoir_weight[14][169],
reservoir_weight[14][170],
reservoir_weight[14][171],
reservoir_weight[14][172],
reservoir_weight[14][173],
reservoir_weight[14][174],
reservoir_weight[14][175],
reservoir_weight[14][176],
reservoir_weight[14][177],
reservoir_weight[14][178],
reservoir_weight[14][179],
reservoir_weight[14][180],
reservoir_weight[14][181],
reservoir_weight[14][182],
reservoir_weight[14][183],
reservoir_weight[14][184],
reservoir_weight[14][185],
reservoir_weight[14][186],
reservoir_weight[14][187],
reservoir_weight[14][188],
reservoir_weight[14][189],
reservoir_weight[14][190],
reservoir_weight[14][191],
reservoir_weight[14][192],
reservoir_weight[14][193],
reservoir_weight[14][194],
reservoir_weight[14][195],
reservoir_weight[14][196],
reservoir_weight[14][197],
reservoir_weight[14][198],
reservoir_weight[14][199]
},
{reservoir_weight[15][0],
reservoir_weight[15][1],
reservoir_weight[15][2],
reservoir_weight[15][3],
reservoir_weight[15][4],
reservoir_weight[15][5],
reservoir_weight[15][6],
reservoir_weight[15][7],
reservoir_weight[15][8],
reservoir_weight[15][9],
reservoir_weight[15][10],
reservoir_weight[15][11],
reservoir_weight[15][12],
reservoir_weight[15][13],
reservoir_weight[15][14],
reservoir_weight[15][15],
reservoir_weight[15][16],
reservoir_weight[15][17],
reservoir_weight[15][18],
reservoir_weight[15][19],
reservoir_weight[15][20],
reservoir_weight[15][21],
reservoir_weight[15][22],
reservoir_weight[15][23],
reservoir_weight[15][24],
reservoir_weight[15][25],
reservoir_weight[15][26],
reservoir_weight[15][27],
reservoir_weight[15][28],
reservoir_weight[15][29],
reservoir_weight[15][30],
reservoir_weight[15][31],
reservoir_weight[15][32],
reservoir_weight[15][33],
reservoir_weight[15][34],
reservoir_weight[15][35],
reservoir_weight[15][36],
reservoir_weight[15][37],
reservoir_weight[15][38],
reservoir_weight[15][39],
reservoir_weight[15][40],
reservoir_weight[15][41],
reservoir_weight[15][42],
reservoir_weight[15][43],
reservoir_weight[15][44],
reservoir_weight[15][45],
reservoir_weight[15][46],
reservoir_weight[15][47],
reservoir_weight[15][48],
reservoir_weight[15][49],
reservoir_weight[15][50],
reservoir_weight[15][51],
reservoir_weight[15][52],
reservoir_weight[15][53],
reservoir_weight[15][54],
reservoir_weight[15][55],
reservoir_weight[15][56],
reservoir_weight[15][57],
reservoir_weight[15][58],
reservoir_weight[15][59],
reservoir_weight[15][60],
reservoir_weight[15][61],
reservoir_weight[15][62],
reservoir_weight[15][63],
reservoir_weight[15][64],
reservoir_weight[15][65],
reservoir_weight[15][66],
reservoir_weight[15][67],
reservoir_weight[15][68],
reservoir_weight[15][69],
reservoir_weight[15][70],
reservoir_weight[15][71],
reservoir_weight[15][72],
reservoir_weight[15][73],
reservoir_weight[15][74],
reservoir_weight[15][75],
reservoir_weight[15][76],
reservoir_weight[15][77],
reservoir_weight[15][78],
reservoir_weight[15][79],
reservoir_weight[15][80],
reservoir_weight[15][81],
reservoir_weight[15][82],
reservoir_weight[15][83],
reservoir_weight[15][84],
reservoir_weight[15][85],
reservoir_weight[15][86],
reservoir_weight[15][87],
reservoir_weight[15][88],
reservoir_weight[15][89],
reservoir_weight[15][90],
reservoir_weight[15][91],
reservoir_weight[15][92],
reservoir_weight[15][93],
reservoir_weight[15][94],
reservoir_weight[15][95],
reservoir_weight[15][96],
reservoir_weight[15][97],
reservoir_weight[15][98],
reservoir_weight[15][99],
reservoir_weight[15][100],
reservoir_weight[15][101],
reservoir_weight[15][102],
reservoir_weight[15][103],
reservoir_weight[15][104],
reservoir_weight[15][105],
reservoir_weight[15][106],
reservoir_weight[15][107],
reservoir_weight[15][108],
reservoir_weight[15][109],
reservoir_weight[15][110],
reservoir_weight[15][111],
reservoir_weight[15][112],
reservoir_weight[15][113],
reservoir_weight[15][114],
reservoir_weight[15][115],
reservoir_weight[15][116],
reservoir_weight[15][117],
reservoir_weight[15][118],
reservoir_weight[15][119],
reservoir_weight[15][120],
reservoir_weight[15][121],
reservoir_weight[15][122],
reservoir_weight[15][123],
reservoir_weight[15][124],
reservoir_weight[15][125],
reservoir_weight[15][126],
reservoir_weight[15][127],
reservoir_weight[15][128],
reservoir_weight[15][129],
reservoir_weight[15][130],
reservoir_weight[15][131],
reservoir_weight[15][132],
reservoir_weight[15][133],
reservoir_weight[15][134],
reservoir_weight[15][135],
reservoir_weight[15][136],
reservoir_weight[15][137],
reservoir_weight[15][138],
reservoir_weight[15][139],
reservoir_weight[15][140],
reservoir_weight[15][141],
reservoir_weight[15][142],
reservoir_weight[15][143],
reservoir_weight[15][144],
reservoir_weight[15][145],
reservoir_weight[15][146],
reservoir_weight[15][147],
reservoir_weight[15][148],
reservoir_weight[15][149],
reservoir_weight[15][150],
reservoir_weight[15][151],
reservoir_weight[15][152],
reservoir_weight[15][153],
reservoir_weight[15][154],
reservoir_weight[15][155],
reservoir_weight[15][156],
reservoir_weight[15][157],
reservoir_weight[15][158],
reservoir_weight[15][159],
reservoir_weight[15][160],
reservoir_weight[15][161],
reservoir_weight[15][162],
reservoir_weight[15][163],
reservoir_weight[15][164],
reservoir_weight[15][165],
reservoir_weight[15][166],
reservoir_weight[15][167],
reservoir_weight[15][168],
reservoir_weight[15][169],
reservoir_weight[15][170],
reservoir_weight[15][171],
reservoir_weight[15][172],
reservoir_weight[15][173],
reservoir_weight[15][174],
reservoir_weight[15][175],
reservoir_weight[15][176],
reservoir_weight[15][177],
reservoir_weight[15][178],
reservoir_weight[15][179],
reservoir_weight[15][180],
reservoir_weight[15][181],
reservoir_weight[15][182],
reservoir_weight[15][183],
reservoir_weight[15][184],
reservoir_weight[15][185],
reservoir_weight[15][186],
reservoir_weight[15][187],
reservoir_weight[15][188],
reservoir_weight[15][189],
reservoir_weight[15][190],
reservoir_weight[15][191],
reservoir_weight[15][192],
reservoir_weight[15][193],
reservoir_weight[15][194],
reservoir_weight[15][195],
reservoir_weight[15][196],
reservoir_weight[15][197],
reservoir_weight[15][198],
reservoir_weight[15][199]
},
{reservoir_weight[16][0],
reservoir_weight[16][1],
reservoir_weight[16][2],
reservoir_weight[16][3],
reservoir_weight[16][4],
reservoir_weight[16][5],
reservoir_weight[16][6],
reservoir_weight[16][7],
reservoir_weight[16][8],
reservoir_weight[16][9],
reservoir_weight[16][10],
reservoir_weight[16][11],
reservoir_weight[16][12],
reservoir_weight[16][13],
reservoir_weight[16][14],
reservoir_weight[16][15],
reservoir_weight[16][16],
reservoir_weight[16][17],
reservoir_weight[16][18],
reservoir_weight[16][19],
reservoir_weight[16][20],
reservoir_weight[16][21],
reservoir_weight[16][22],
reservoir_weight[16][23],
reservoir_weight[16][24],
reservoir_weight[16][25],
reservoir_weight[16][26],
reservoir_weight[16][27],
reservoir_weight[16][28],
reservoir_weight[16][29],
reservoir_weight[16][30],
reservoir_weight[16][31],
reservoir_weight[16][32],
reservoir_weight[16][33],
reservoir_weight[16][34],
reservoir_weight[16][35],
reservoir_weight[16][36],
reservoir_weight[16][37],
reservoir_weight[16][38],
reservoir_weight[16][39],
reservoir_weight[16][40],
reservoir_weight[16][41],
reservoir_weight[16][42],
reservoir_weight[16][43],
reservoir_weight[16][44],
reservoir_weight[16][45],
reservoir_weight[16][46],
reservoir_weight[16][47],
reservoir_weight[16][48],
reservoir_weight[16][49],
reservoir_weight[16][50],
reservoir_weight[16][51],
reservoir_weight[16][52],
reservoir_weight[16][53],
reservoir_weight[16][54],
reservoir_weight[16][55],
reservoir_weight[16][56],
reservoir_weight[16][57],
reservoir_weight[16][58],
reservoir_weight[16][59],
reservoir_weight[16][60],
reservoir_weight[16][61],
reservoir_weight[16][62],
reservoir_weight[16][63],
reservoir_weight[16][64],
reservoir_weight[16][65],
reservoir_weight[16][66],
reservoir_weight[16][67],
reservoir_weight[16][68],
reservoir_weight[16][69],
reservoir_weight[16][70],
reservoir_weight[16][71],
reservoir_weight[16][72],
reservoir_weight[16][73],
reservoir_weight[16][74],
reservoir_weight[16][75],
reservoir_weight[16][76],
reservoir_weight[16][77],
reservoir_weight[16][78],
reservoir_weight[16][79],
reservoir_weight[16][80],
reservoir_weight[16][81],
reservoir_weight[16][82],
reservoir_weight[16][83],
reservoir_weight[16][84],
reservoir_weight[16][85],
reservoir_weight[16][86],
reservoir_weight[16][87],
reservoir_weight[16][88],
reservoir_weight[16][89],
reservoir_weight[16][90],
reservoir_weight[16][91],
reservoir_weight[16][92],
reservoir_weight[16][93],
reservoir_weight[16][94],
reservoir_weight[16][95],
reservoir_weight[16][96],
reservoir_weight[16][97],
reservoir_weight[16][98],
reservoir_weight[16][99],
reservoir_weight[16][100],
reservoir_weight[16][101],
reservoir_weight[16][102],
reservoir_weight[16][103],
reservoir_weight[16][104],
reservoir_weight[16][105],
reservoir_weight[16][106],
reservoir_weight[16][107],
reservoir_weight[16][108],
reservoir_weight[16][109],
reservoir_weight[16][110],
reservoir_weight[16][111],
reservoir_weight[16][112],
reservoir_weight[16][113],
reservoir_weight[16][114],
reservoir_weight[16][115],
reservoir_weight[16][116],
reservoir_weight[16][117],
reservoir_weight[16][118],
reservoir_weight[16][119],
reservoir_weight[16][120],
reservoir_weight[16][121],
reservoir_weight[16][122],
reservoir_weight[16][123],
reservoir_weight[16][124],
reservoir_weight[16][125],
reservoir_weight[16][126],
reservoir_weight[16][127],
reservoir_weight[16][128],
reservoir_weight[16][129],
reservoir_weight[16][130],
reservoir_weight[16][131],
reservoir_weight[16][132],
reservoir_weight[16][133],
reservoir_weight[16][134],
reservoir_weight[16][135],
reservoir_weight[16][136],
reservoir_weight[16][137],
reservoir_weight[16][138],
reservoir_weight[16][139],
reservoir_weight[16][140],
reservoir_weight[16][141],
reservoir_weight[16][142],
reservoir_weight[16][143],
reservoir_weight[16][144],
reservoir_weight[16][145],
reservoir_weight[16][146],
reservoir_weight[16][147],
reservoir_weight[16][148],
reservoir_weight[16][149],
reservoir_weight[16][150],
reservoir_weight[16][151],
reservoir_weight[16][152],
reservoir_weight[16][153],
reservoir_weight[16][154],
reservoir_weight[16][155],
reservoir_weight[16][156],
reservoir_weight[16][157],
reservoir_weight[16][158],
reservoir_weight[16][159],
reservoir_weight[16][160],
reservoir_weight[16][161],
reservoir_weight[16][162],
reservoir_weight[16][163],
reservoir_weight[16][164],
reservoir_weight[16][165],
reservoir_weight[16][166],
reservoir_weight[16][167],
reservoir_weight[16][168],
reservoir_weight[16][169],
reservoir_weight[16][170],
reservoir_weight[16][171],
reservoir_weight[16][172],
reservoir_weight[16][173],
reservoir_weight[16][174],
reservoir_weight[16][175],
reservoir_weight[16][176],
reservoir_weight[16][177],
reservoir_weight[16][178],
reservoir_weight[16][179],
reservoir_weight[16][180],
reservoir_weight[16][181],
reservoir_weight[16][182],
reservoir_weight[16][183],
reservoir_weight[16][184],
reservoir_weight[16][185],
reservoir_weight[16][186],
reservoir_weight[16][187],
reservoir_weight[16][188],
reservoir_weight[16][189],
reservoir_weight[16][190],
reservoir_weight[16][191],
reservoir_weight[16][192],
reservoir_weight[16][193],
reservoir_weight[16][194],
reservoir_weight[16][195],
reservoir_weight[16][196],
reservoir_weight[16][197],
reservoir_weight[16][198],
reservoir_weight[16][199]
},
{reservoir_weight[17][0],
reservoir_weight[17][1],
reservoir_weight[17][2],
reservoir_weight[17][3],
reservoir_weight[17][4],
reservoir_weight[17][5],
reservoir_weight[17][6],
reservoir_weight[17][7],
reservoir_weight[17][8],
reservoir_weight[17][9],
reservoir_weight[17][10],
reservoir_weight[17][11],
reservoir_weight[17][12],
reservoir_weight[17][13],
reservoir_weight[17][14],
reservoir_weight[17][15],
reservoir_weight[17][16],
reservoir_weight[17][17],
reservoir_weight[17][18],
reservoir_weight[17][19],
reservoir_weight[17][20],
reservoir_weight[17][21],
reservoir_weight[17][22],
reservoir_weight[17][23],
reservoir_weight[17][24],
reservoir_weight[17][25],
reservoir_weight[17][26],
reservoir_weight[17][27],
reservoir_weight[17][28],
reservoir_weight[17][29],
reservoir_weight[17][30],
reservoir_weight[17][31],
reservoir_weight[17][32],
reservoir_weight[17][33],
reservoir_weight[17][34],
reservoir_weight[17][35],
reservoir_weight[17][36],
reservoir_weight[17][37],
reservoir_weight[17][38],
reservoir_weight[17][39],
reservoir_weight[17][40],
reservoir_weight[17][41],
reservoir_weight[17][42],
reservoir_weight[17][43],
reservoir_weight[17][44],
reservoir_weight[17][45],
reservoir_weight[17][46],
reservoir_weight[17][47],
reservoir_weight[17][48],
reservoir_weight[17][49],
reservoir_weight[17][50],
reservoir_weight[17][51],
reservoir_weight[17][52],
reservoir_weight[17][53],
reservoir_weight[17][54],
reservoir_weight[17][55],
reservoir_weight[17][56],
reservoir_weight[17][57],
reservoir_weight[17][58],
reservoir_weight[17][59],
reservoir_weight[17][60],
reservoir_weight[17][61],
reservoir_weight[17][62],
reservoir_weight[17][63],
reservoir_weight[17][64],
reservoir_weight[17][65],
reservoir_weight[17][66],
reservoir_weight[17][67],
reservoir_weight[17][68],
reservoir_weight[17][69],
reservoir_weight[17][70],
reservoir_weight[17][71],
reservoir_weight[17][72],
reservoir_weight[17][73],
reservoir_weight[17][74],
reservoir_weight[17][75],
reservoir_weight[17][76],
reservoir_weight[17][77],
reservoir_weight[17][78],
reservoir_weight[17][79],
reservoir_weight[17][80],
reservoir_weight[17][81],
reservoir_weight[17][82],
reservoir_weight[17][83],
reservoir_weight[17][84],
reservoir_weight[17][85],
reservoir_weight[17][86],
reservoir_weight[17][87],
reservoir_weight[17][88],
reservoir_weight[17][89],
reservoir_weight[17][90],
reservoir_weight[17][91],
reservoir_weight[17][92],
reservoir_weight[17][93],
reservoir_weight[17][94],
reservoir_weight[17][95],
reservoir_weight[17][96],
reservoir_weight[17][97],
reservoir_weight[17][98],
reservoir_weight[17][99],
reservoir_weight[17][100],
reservoir_weight[17][101],
reservoir_weight[17][102],
reservoir_weight[17][103],
reservoir_weight[17][104],
reservoir_weight[17][105],
reservoir_weight[17][106],
reservoir_weight[17][107],
reservoir_weight[17][108],
reservoir_weight[17][109],
reservoir_weight[17][110],
reservoir_weight[17][111],
reservoir_weight[17][112],
reservoir_weight[17][113],
reservoir_weight[17][114],
reservoir_weight[17][115],
reservoir_weight[17][116],
reservoir_weight[17][117],
reservoir_weight[17][118],
reservoir_weight[17][119],
reservoir_weight[17][120],
reservoir_weight[17][121],
reservoir_weight[17][122],
reservoir_weight[17][123],
reservoir_weight[17][124],
reservoir_weight[17][125],
reservoir_weight[17][126],
reservoir_weight[17][127],
reservoir_weight[17][128],
reservoir_weight[17][129],
reservoir_weight[17][130],
reservoir_weight[17][131],
reservoir_weight[17][132],
reservoir_weight[17][133],
reservoir_weight[17][134],
reservoir_weight[17][135],
reservoir_weight[17][136],
reservoir_weight[17][137],
reservoir_weight[17][138],
reservoir_weight[17][139],
reservoir_weight[17][140],
reservoir_weight[17][141],
reservoir_weight[17][142],
reservoir_weight[17][143],
reservoir_weight[17][144],
reservoir_weight[17][145],
reservoir_weight[17][146],
reservoir_weight[17][147],
reservoir_weight[17][148],
reservoir_weight[17][149],
reservoir_weight[17][150],
reservoir_weight[17][151],
reservoir_weight[17][152],
reservoir_weight[17][153],
reservoir_weight[17][154],
reservoir_weight[17][155],
reservoir_weight[17][156],
reservoir_weight[17][157],
reservoir_weight[17][158],
reservoir_weight[17][159],
reservoir_weight[17][160],
reservoir_weight[17][161],
reservoir_weight[17][162],
reservoir_weight[17][163],
reservoir_weight[17][164],
reservoir_weight[17][165],
reservoir_weight[17][166],
reservoir_weight[17][167],
reservoir_weight[17][168],
reservoir_weight[17][169],
reservoir_weight[17][170],
reservoir_weight[17][171],
reservoir_weight[17][172],
reservoir_weight[17][173],
reservoir_weight[17][174],
reservoir_weight[17][175],
reservoir_weight[17][176],
reservoir_weight[17][177],
reservoir_weight[17][178],
reservoir_weight[17][179],
reservoir_weight[17][180],
reservoir_weight[17][181],
reservoir_weight[17][182],
reservoir_weight[17][183],
reservoir_weight[17][184],
reservoir_weight[17][185],
reservoir_weight[17][186],
reservoir_weight[17][187],
reservoir_weight[17][188],
reservoir_weight[17][189],
reservoir_weight[17][190],
reservoir_weight[17][191],
reservoir_weight[17][192],
reservoir_weight[17][193],
reservoir_weight[17][194],
reservoir_weight[17][195],
reservoir_weight[17][196],
reservoir_weight[17][197],
reservoir_weight[17][198],
reservoir_weight[17][199]
},
{reservoir_weight[18][0],
reservoir_weight[18][1],
reservoir_weight[18][2],
reservoir_weight[18][3],
reservoir_weight[18][4],
reservoir_weight[18][5],
reservoir_weight[18][6],
reservoir_weight[18][7],
reservoir_weight[18][8],
reservoir_weight[18][9],
reservoir_weight[18][10],
reservoir_weight[18][11],
reservoir_weight[18][12],
reservoir_weight[18][13],
reservoir_weight[18][14],
reservoir_weight[18][15],
reservoir_weight[18][16],
reservoir_weight[18][17],
reservoir_weight[18][18],
reservoir_weight[18][19],
reservoir_weight[18][20],
reservoir_weight[18][21],
reservoir_weight[18][22],
reservoir_weight[18][23],
reservoir_weight[18][24],
reservoir_weight[18][25],
reservoir_weight[18][26],
reservoir_weight[18][27],
reservoir_weight[18][28],
reservoir_weight[18][29],
reservoir_weight[18][30],
reservoir_weight[18][31],
reservoir_weight[18][32],
reservoir_weight[18][33],
reservoir_weight[18][34],
reservoir_weight[18][35],
reservoir_weight[18][36],
reservoir_weight[18][37],
reservoir_weight[18][38],
reservoir_weight[18][39],
reservoir_weight[18][40],
reservoir_weight[18][41],
reservoir_weight[18][42],
reservoir_weight[18][43],
reservoir_weight[18][44],
reservoir_weight[18][45],
reservoir_weight[18][46],
reservoir_weight[18][47],
reservoir_weight[18][48],
reservoir_weight[18][49],
reservoir_weight[18][50],
reservoir_weight[18][51],
reservoir_weight[18][52],
reservoir_weight[18][53],
reservoir_weight[18][54],
reservoir_weight[18][55],
reservoir_weight[18][56],
reservoir_weight[18][57],
reservoir_weight[18][58],
reservoir_weight[18][59],
reservoir_weight[18][60],
reservoir_weight[18][61],
reservoir_weight[18][62],
reservoir_weight[18][63],
reservoir_weight[18][64],
reservoir_weight[18][65],
reservoir_weight[18][66],
reservoir_weight[18][67],
reservoir_weight[18][68],
reservoir_weight[18][69],
reservoir_weight[18][70],
reservoir_weight[18][71],
reservoir_weight[18][72],
reservoir_weight[18][73],
reservoir_weight[18][74],
reservoir_weight[18][75],
reservoir_weight[18][76],
reservoir_weight[18][77],
reservoir_weight[18][78],
reservoir_weight[18][79],
reservoir_weight[18][80],
reservoir_weight[18][81],
reservoir_weight[18][82],
reservoir_weight[18][83],
reservoir_weight[18][84],
reservoir_weight[18][85],
reservoir_weight[18][86],
reservoir_weight[18][87],
reservoir_weight[18][88],
reservoir_weight[18][89],
reservoir_weight[18][90],
reservoir_weight[18][91],
reservoir_weight[18][92],
reservoir_weight[18][93],
reservoir_weight[18][94],
reservoir_weight[18][95],
reservoir_weight[18][96],
reservoir_weight[18][97],
reservoir_weight[18][98],
reservoir_weight[18][99],
reservoir_weight[18][100],
reservoir_weight[18][101],
reservoir_weight[18][102],
reservoir_weight[18][103],
reservoir_weight[18][104],
reservoir_weight[18][105],
reservoir_weight[18][106],
reservoir_weight[18][107],
reservoir_weight[18][108],
reservoir_weight[18][109],
reservoir_weight[18][110],
reservoir_weight[18][111],
reservoir_weight[18][112],
reservoir_weight[18][113],
reservoir_weight[18][114],
reservoir_weight[18][115],
reservoir_weight[18][116],
reservoir_weight[18][117],
reservoir_weight[18][118],
reservoir_weight[18][119],
reservoir_weight[18][120],
reservoir_weight[18][121],
reservoir_weight[18][122],
reservoir_weight[18][123],
reservoir_weight[18][124],
reservoir_weight[18][125],
reservoir_weight[18][126],
reservoir_weight[18][127],
reservoir_weight[18][128],
reservoir_weight[18][129],
reservoir_weight[18][130],
reservoir_weight[18][131],
reservoir_weight[18][132],
reservoir_weight[18][133],
reservoir_weight[18][134],
reservoir_weight[18][135],
reservoir_weight[18][136],
reservoir_weight[18][137],
reservoir_weight[18][138],
reservoir_weight[18][139],
reservoir_weight[18][140],
reservoir_weight[18][141],
reservoir_weight[18][142],
reservoir_weight[18][143],
reservoir_weight[18][144],
reservoir_weight[18][145],
reservoir_weight[18][146],
reservoir_weight[18][147],
reservoir_weight[18][148],
reservoir_weight[18][149],
reservoir_weight[18][150],
reservoir_weight[18][151],
reservoir_weight[18][152],
reservoir_weight[18][153],
reservoir_weight[18][154],
reservoir_weight[18][155],
reservoir_weight[18][156],
reservoir_weight[18][157],
reservoir_weight[18][158],
reservoir_weight[18][159],
reservoir_weight[18][160],
reservoir_weight[18][161],
reservoir_weight[18][162],
reservoir_weight[18][163],
reservoir_weight[18][164],
reservoir_weight[18][165],
reservoir_weight[18][166],
reservoir_weight[18][167],
reservoir_weight[18][168],
reservoir_weight[18][169],
reservoir_weight[18][170],
reservoir_weight[18][171],
reservoir_weight[18][172],
reservoir_weight[18][173],
reservoir_weight[18][174],
reservoir_weight[18][175],
reservoir_weight[18][176],
reservoir_weight[18][177],
reservoir_weight[18][178],
reservoir_weight[18][179],
reservoir_weight[18][180],
reservoir_weight[18][181],
reservoir_weight[18][182],
reservoir_weight[18][183],
reservoir_weight[18][184],
reservoir_weight[18][185],
reservoir_weight[18][186],
reservoir_weight[18][187],
reservoir_weight[18][188],
reservoir_weight[18][189],
reservoir_weight[18][190],
reservoir_weight[18][191],
reservoir_weight[18][192],
reservoir_weight[18][193],
reservoir_weight[18][194],
reservoir_weight[18][195],
reservoir_weight[18][196],
reservoir_weight[18][197],
reservoir_weight[18][198],
reservoir_weight[18][199]
},
{reservoir_weight[19][0],
reservoir_weight[19][1],
reservoir_weight[19][2],
reservoir_weight[19][3],
reservoir_weight[19][4],
reservoir_weight[19][5],
reservoir_weight[19][6],
reservoir_weight[19][7],
reservoir_weight[19][8],
reservoir_weight[19][9],
reservoir_weight[19][10],
reservoir_weight[19][11],
reservoir_weight[19][12],
reservoir_weight[19][13],
reservoir_weight[19][14],
reservoir_weight[19][15],
reservoir_weight[19][16],
reservoir_weight[19][17],
reservoir_weight[19][18],
reservoir_weight[19][19],
reservoir_weight[19][20],
reservoir_weight[19][21],
reservoir_weight[19][22],
reservoir_weight[19][23],
reservoir_weight[19][24],
reservoir_weight[19][25],
reservoir_weight[19][26],
reservoir_weight[19][27],
reservoir_weight[19][28],
reservoir_weight[19][29],
reservoir_weight[19][30],
reservoir_weight[19][31],
reservoir_weight[19][32],
reservoir_weight[19][33],
reservoir_weight[19][34],
reservoir_weight[19][35],
reservoir_weight[19][36],
reservoir_weight[19][37],
reservoir_weight[19][38],
reservoir_weight[19][39],
reservoir_weight[19][40],
reservoir_weight[19][41],
reservoir_weight[19][42],
reservoir_weight[19][43],
reservoir_weight[19][44],
reservoir_weight[19][45],
reservoir_weight[19][46],
reservoir_weight[19][47],
reservoir_weight[19][48],
reservoir_weight[19][49],
reservoir_weight[19][50],
reservoir_weight[19][51],
reservoir_weight[19][52],
reservoir_weight[19][53],
reservoir_weight[19][54],
reservoir_weight[19][55],
reservoir_weight[19][56],
reservoir_weight[19][57],
reservoir_weight[19][58],
reservoir_weight[19][59],
reservoir_weight[19][60],
reservoir_weight[19][61],
reservoir_weight[19][62],
reservoir_weight[19][63],
reservoir_weight[19][64],
reservoir_weight[19][65],
reservoir_weight[19][66],
reservoir_weight[19][67],
reservoir_weight[19][68],
reservoir_weight[19][69],
reservoir_weight[19][70],
reservoir_weight[19][71],
reservoir_weight[19][72],
reservoir_weight[19][73],
reservoir_weight[19][74],
reservoir_weight[19][75],
reservoir_weight[19][76],
reservoir_weight[19][77],
reservoir_weight[19][78],
reservoir_weight[19][79],
reservoir_weight[19][80],
reservoir_weight[19][81],
reservoir_weight[19][82],
reservoir_weight[19][83],
reservoir_weight[19][84],
reservoir_weight[19][85],
reservoir_weight[19][86],
reservoir_weight[19][87],
reservoir_weight[19][88],
reservoir_weight[19][89],
reservoir_weight[19][90],
reservoir_weight[19][91],
reservoir_weight[19][92],
reservoir_weight[19][93],
reservoir_weight[19][94],
reservoir_weight[19][95],
reservoir_weight[19][96],
reservoir_weight[19][97],
reservoir_weight[19][98],
reservoir_weight[19][99],
reservoir_weight[19][100],
reservoir_weight[19][101],
reservoir_weight[19][102],
reservoir_weight[19][103],
reservoir_weight[19][104],
reservoir_weight[19][105],
reservoir_weight[19][106],
reservoir_weight[19][107],
reservoir_weight[19][108],
reservoir_weight[19][109],
reservoir_weight[19][110],
reservoir_weight[19][111],
reservoir_weight[19][112],
reservoir_weight[19][113],
reservoir_weight[19][114],
reservoir_weight[19][115],
reservoir_weight[19][116],
reservoir_weight[19][117],
reservoir_weight[19][118],
reservoir_weight[19][119],
reservoir_weight[19][120],
reservoir_weight[19][121],
reservoir_weight[19][122],
reservoir_weight[19][123],
reservoir_weight[19][124],
reservoir_weight[19][125],
reservoir_weight[19][126],
reservoir_weight[19][127],
reservoir_weight[19][128],
reservoir_weight[19][129],
reservoir_weight[19][130],
reservoir_weight[19][131],
reservoir_weight[19][132],
reservoir_weight[19][133],
reservoir_weight[19][134],
reservoir_weight[19][135],
reservoir_weight[19][136],
reservoir_weight[19][137],
reservoir_weight[19][138],
reservoir_weight[19][139],
reservoir_weight[19][140],
reservoir_weight[19][141],
reservoir_weight[19][142],
reservoir_weight[19][143],
reservoir_weight[19][144],
reservoir_weight[19][145],
reservoir_weight[19][146],
reservoir_weight[19][147],
reservoir_weight[19][148],
reservoir_weight[19][149],
reservoir_weight[19][150],
reservoir_weight[19][151],
reservoir_weight[19][152],
reservoir_weight[19][153],
reservoir_weight[19][154],
reservoir_weight[19][155],
reservoir_weight[19][156],
reservoir_weight[19][157],
reservoir_weight[19][158],
reservoir_weight[19][159],
reservoir_weight[19][160],
reservoir_weight[19][161],
reservoir_weight[19][162],
reservoir_weight[19][163],
reservoir_weight[19][164],
reservoir_weight[19][165],
reservoir_weight[19][166],
reservoir_weight[19][167],
reservoir_weight[19][168],
reservoir_weight[19][169],
reservoir_weight[19][170],
reservoir_weight[19][171],
reservoir_weight[19][172],
reservoir_weight[19][173],
reservoir_weight[19][174],
reservoir_weight[19][175],
reservoir_weight[19][176],
reservoir_weight[19][177],
reservoir_weight[19][178],
reservoir_weight[19][179],
reservoir_weight[19][180],
reservoir_weight[19][181],
reservoir_weight[19][182],
reservoir_weight[19][183],
reservoir_weight[19][184],
reservoir_weight[19][185],
reservoir_weight[19][186],
reservoir_weight[19][187],
reservoir_weight[19][188],
reservoir_weight[19][189],
reservoir_weight[19][190],
reservoir_weight[19][191],
reservoir_weight[19][192],
reservoir_weight[19][193],
reservoir_weight[19][194],
reservoir_weight[19][195],
reservoir_weight[19][196],
reservoir_weight[19][197],
reservoir_weight[19][198],
reservoir_weight[19][199]
},
{reservoir_weight[20][0],
reservoir_weight[20][1],
reservoir_weight[20][2],
reservoir_weight[20][3],
reservoir_weight[20][4],
reservoir_weight[20][5],
reservoir_weight[20][6],
reservoir_weight[20][7],
reservoir_weight[20][8],
reservoir_weight[20][9],
reservoir_weight[20][10],
reservoir_weight[20][11],
reservoir_weight[20][12],
reservoir_weight[20][13],
reservoir_weight[20][14],
reservoir_weight[20][15],
reservoir_weight[20][16],
reservoir_weight[20][17],
reservoir_weight[20][18],
reservoir_weight[20][19],
reservoir_weight[20][20],
reservoir_weight[20][21],
reservoir_weight[20][22],
reservoir_weight[20][23],
reservoir_weight[20][24],
reservoir_weight[20][25],
reservoir_weight[20][26],
reservoir_weight[20][27],
reservoir_weight[20][28],
reservoir_weight[20][29],
reservoir_weight[20][30],
reservoir_weight[20][31],
reservoir_weight[20][32],
reservoir_weight[20][33],
reservoir_weight[20][34],
reservoir_weight[20][35],
reservoir_weight[20][36],
reservoir_weight[20][37],
reservoir_weight[20][38],
reservoir_weight[20][39],
reservoir_weight[20][40],
reservoir_weight[20][41],
reservoir_weight[20][42],
reservoir_weight[20][43],
reservoir_weight[20][44],
reservoir_weight[20][45],
reservoir_weight[20][46],
reservoir_weight[20][47],
reservoir_weight[20][48],
reservoir_weight[20][49],
reservoir_weight[20][50],
reservoir_weight[20][51],
reservoir_weight[20][52],
reservoir_weight[20][53],
reservoir_weight[20][54],
reservoir_weight[20][55],
reservoir_weight[20][56],
reservoir_weight[20][57],
reservoir_weight[20][58],
reservoir_weight[20][59],
reservoir_weight[20][60],
reservoir_weight[20][61],
reservoir_weight[20][62],
reservoir_weight[20][63],
reservoir_weight[20][64],
reservoir_weight[20][65],
reservoir_weight[20][66],
reservoir_weight[20][67],
reservoir_weight[20][68],
reservoir_weight[20][69],
reservoir_weight[20][70],
reservoir_weight[20][71],
reservoir_weight[20][72],
reservoir_weight[20][73],
reservoir_weight[20][74],
reservoir_weight[20][75],
reservoir_weight[20][76],
reservoir_weight[20][77],
reservoir_weight[20][78],
reservoir_weight[20][79],
reservoir_weight[20][80],
reservoir_weight[20][81],
reservoir_weight[20][82],
reservoir_weight[20][83],
reservoir_weight[20][84],
reservoir_weight[20][85],
reservoir_weight[20][86],
reservoir_weight[20][87],
reservoir_weight[20][88],
reservoir_weight[20][89],
reservoir_weight[20][90],
reservoir_weight[20][91],
reservoir_weight[20][92],
reservoir_weight[20][93],
reservoir_weight[20][94],
reservoir_weight[20][95],
reservoir_weight[20][96],
reservoir_weight[20][97],
reservoir_weight[20][98],
reservoir_weight[20][99],
reservoir_weight[20][100],
reservoir_weight[20][101],
reservoir_weight[20][102],
reservoir_weight[20][103],
reservoir_weight[20][104],
reservoir_weight[20][105],
reservoir_weight[20][106],
reservoir_weight[20][107],
reservoir_weight[20][108],
reservoir_weight[20][109],
reservoir_weight[20][110],
reservoir_weight[20][111],
reservoir_weight[20][112],
reservoir_weight[20][113],
reservoir_weight[20][114],
reservoir_weight[20][115],
reservoir_weight[20][116],
reservoir_weight[20][117],
reservoir_weight[20][118],
reservoir_weight[20][119],
reservoir_weight[20][120],
reservoir_weight[20][121],
reservoir_weight[20][122],
reservoir_weight[20][123],
reservoir_weight[20][124],
reservoir_weight[20][125],
reservoir_weight[20][126],
reservoir_weight[20][127],
reservoir_weight[20][128],
reservoir_weight[20][129],
reservoir_weight[20][130],
reservoir_weight[20][131],
reservoir_weight[20][132],
reservoir_weight[20][133],
reservoir_weight[20][134],
reservoir_weight[20][135],
reservoir_weight[20][136],
reservoir_weight[20][137],
reservoir_weight[20][138],
reservoir_weight[20][139],
reservoir_weight[20][140],
reservoir_weight[20][141],
reservoir_weight[20][142],
reservoir_weight[20][143],
reservoir_weight[20][144],
reservoir_weight[20][145],
reservoir_weight[20][146],
reservoir_weight[20][147],
reservoir_weight[20][148],
reservoir_weight[20][149],
reservoir_weight[20][150],
reservoir_weight[20][151],
reservoir_weight[20][152],
reservoir_weight[20][153],
reservoir_weight[20][154],
reservoir_weight[20][155],
reservoir_weight[20][156],
reservoir_weight[20][157],
reservoir_weight[20][158],
reservoir_weight[20][159],
reservoir_weight[20][160],
reservoir_weight[20][161],
reservoir_weight[20][162],
reservoir_weight[20][163],
reservoir_weight[20][164],
reservoir_weight[20][165],
reservoir_weight[20][166],
reservoir_weight[20][167],
reservoir_weight[20][168],
reservoir_weight[20][169],
reservoir_weight[20][170],
reservoir_weight[20][171],
reservoir_weight[20][172],
reservoir_weight[20][173],
reservoir_weight[20][174],
reservoir_weight[20][175],
reservoir_weight[20][176],
reservoir_weight[20][177],
reservoir_weight[20][178],
reservoir_weight[20][179],
reservoir_weight[20][180],
reservoir_weight[20][181],
reservoir_weight[20][182],
reservoir_weight[20][183],
reservoir_weight[20][184],
reservoir_weight[20][185],
reservoir_weight[20][186],
reservoir_weight[20][187],
reservoir_weight[20][188],
reservoir_weight[20][189],
reservoir_weight[20][190],
reservoir_weight[20][191],
reservoir_weight[20][192],
reservoir_weight[20][193],
reservoir_weight[20][194],
reservoir_weight[20][195],
reservoir_weight[20][196],
reservoir_weight[20][197],
reservoir_weight[20][198],
reservoir_weight[20][199]
},
{reservoir_weight[21][0],
reservoir_weight[21][1],
reservoir_weight[21][2],
reservoir_weight[21][3],
reservoir_weight[21][4],
reservoir_weight[21][5],
reservoir_weight[21][6],
reservoir_weight[21][7],
reservoir_weight[21][8],
reservoir_weight[21][9],
reservoir_weight[21][10],
reservoir_weight[21][11],
reservoir_weight[21][12],
reservoir_weight[21][13],
reservoir_weight[21][14],
reservoir_weight[21][15],
reservoir_weight[21][16],
reservoir_weight[21][17],
reservoir_weight[21][18],
reservoir_weight[21][19],
reservoir_weight[21][20],
reservoir_weight[21][21],
reservoir_weight[21][22],
reservoir_weight[21][23],
reservoir_weight[21][24],
reservoir_weight[21][25],
reservoir_weight[21][26],
reservoir_weight[21][27],
reservoir_weight[21][28],
reservoir_weight[21][29],
reservoir_weight[21][30],
reservoir_weight[21][31],
reservoir_weight[21][32],
reservoir_weight[21][33],
reservoir_weight[21][34],
reservoir_weight[21][35],
reservoir_weight[21][36],
reservoir_weight[21][37],
reservoir_weight[21][38],
reservoir_weight[21][39],
reservoir_weight[21][40],
reservoir_weight[21][41],
reservoir_weight[21][42],
reservoir_weight[21][43],
reservoir_weight[21][44],
reservoir_weight[21][45],
reservoir_weight[21][46],
reservoir_weight[21][47],
reservoir_weight[21][48],
reservoir_weight[21][49],
reservoir_weight[21][50],
reservoir_weight[21][51],
reservoir_weight[21][52],
reservoir_weight[21][53],
reservoir_weight[21][54],
reservoir_weight[21][55],
reservoir_weight[21][56],
reservoir_weight[21][57],
reservoir_weight[21][58],
reservoir_weight[21][59],
reservoir_weight[21][60],
reservoir_weight[21][61],
reservoir_weight[21][62],
reservoir_weight[21][63],
reservoir_weight[21][64],
reservoir_weight[21][65],
reservoir_weight[21][66],
reservoir_weight[21][67],
reservoir_weight[21][68],
reservoir_weight[21][69],
reservoir_weight[21][70],
reservoir_weight[21][71],
reservoir_weight[21][72],
reservoir_weight[21][73],
reservoir_weight[21][74],
reservoir_weight[21][75],
reservoir_weight[21][76],
reservoir_weight[21][77],
reservoir_weight[21][78],
reservoir_weight[21][79],
reservoir_weight[21][80],
reservoir_weight[21][81],
reservoir_weight[21][82],
reservoir_weight[21][83],
reservoir_weight[21][84],
reservoir_weight[21][85],
reservoir_weight[21][86],
reservoir_weight[21][87],
reservoir_weight[21][88],
reservoir_weight[21][89],
reservoir_weight[21][90],
reservoir_weight[21][91],
reservoir_weight[21][92],
reservoir_weight[21][93],
reservoir_weight[21][94],
reservoir_weight[21][95],
reservoir_weight[21][96],
reservoir_weight[21][97],
reservoir_weight[21][98],
reservoir_weight[21][99],
reservoir_weight[21][100],
reservoir_weight[21][101],
reservoir_weight[21][102],
reservoir_weight[21][103],
reservoir_weight[21][104],
reservoir_weight[21][105],
reservoir_weight[21][106],
reservoir_weight[21][107],
reservoir_weight[21][108],
reservoir_weight[21][109],
reservoir_weight[21][110],
reservoir_weight[21][111],
reservoir_weight[21][112],
reservoir_weight[21][113],
reservoir_weight[21][114],
reservoir_weight[21][115],
reservoir_weight[21][116],
reservoir_weight[21][117],
reservoir_weight[21][118],
reservoir_weight[21][119],
reservoir_weight[21][120],
reservoir_weight[21][121],
reservoir_weight[21][122],
reservoir_weight[21][123],
reservoir_weight[21][124],
reservoir_weight[21][125],
reservoir_weight[21][126],
reservoir_weight[21][127],
reservoir_weight[21][128],
reservoir_weight[21][129],
reservoir_weight[21][130],
reservoir_weight[21][131],
reservoir_weight[21][132],
reservoir_weight[21][133],
reservoir_weight[21][134],
reservoir_weight[21][135],
reservoir_weight[21][136],
reservoir_weight[21][137],
reservoir_weight[21][138],
reservoir_weight[21][139],
reservoir_weight[21][140],
reservoir_weight[21][141],
reservoir_weight[21][142],
reservoir_weight[21][143],
reservoir_weight[21][144],
reservoir_weight[21][145],
reservoir_weight[21][146],
reservoir_weight[21][147],
reservoir_weight[21][148],
reservoir_weight[21][149],
reservoir_weight[21][150],
reservoir_weight[21][151],
reservoir_weight[21][152],
reservoir_weight[21][153],
reservoir_weight[21][154],
reservoir_weight[21][155],
reservoir_weight[21][156],
reservoir_weight[21][157],
reservoir_weight[21][158],
reservoir_weight[21][159],
reservoir_weight[21][160],
reservoir_weight[21][161],
reservoir_weight[21][162],
reservoir_weight[21][163],
reservoir_weight[21][164],
reservoir_weight[21][165],
reservoir_weight[21][166],
reservoir_weight[21][167],
reservoir_weight[21][168],
reservoir_weight[21][169],
reservoir_weight[21][170],
reservoir_weight[21][171],
reservoir_weight[21][172],
reservoir_weight[21][173],
reservoir_weight[21][174],
reservoir_weight[21][175],
reservoir_weight[21][176],
reservoir_weight[21][177],
reservoir_weight[21][178],
reservoir_weight[21][179],
reservoir_weight[21][180],
reservoir_weight[21][181],
reservoir_weight[21][182],
reservoir_weight[21][183],
reservoir_weight[21][184],
reservoir_weight[21][185],
reservoir_weight[21][186],
reservoir_weight[21][187],
reservoir_weight[21][188],
reservoir_weight[21][189],
reservoir_weight[21][190],
reservoir_weight[21][191],
reservoir_weight[21][192],
reservoir_weight[21][193],
reservoir_weight[21][194],
reservoir_weight[21][195],
reservoir_weight[21][196],
reservoir_weight[21][197],
reservoir_weight[21][198],
reservoir_weight[21][199]
},
{reservoir_weight[22][0],
reservoir_weight[22][1],
reservoir_weight[22][2],
reservoir_weight[22][3],
reservoir_weight[22][4],
reservoir_weight[22][5],
reservoir_weight[22][6],
reservoir_weight[22][7],
reservoir_weight[22][8],
reservoir_weight[22][9],
reservoir_weight[22][10],
reservoir_weight[22][11],
reservoir_weight[22][12],
reservoir_weight[22][13],
reservoir_weight[22][14],
reservoir_weight[22][15],
reservoir_weight[22][16],
reservoir_weight[22][17],
reservoir_weight[22][18],
reservoir_weight[22][19],
reservoir_weight[22][20],
reservoir_weight[22][21],
reservoir_weight[22][22],
reservoir_weight[22][23],
reservoir_weight[22][24],
reservoir_weight[22][25],
reservoir_weight[22][26],
reservoir_weight[22][27],
reservoir_weight[22][28],
reservoir_weight[22][29],
reservoir_weight[22][30],
reservoir_weight[22][31],
reservoir_weight[22][32],
reservoir_weight[22][33],
reservoir_weight[22][34],
reservoir_weight[22][35],
reservoir_weight[22][36],
reservoir_weight[22][37],
reservoir_weight[22][38],
reservoir_weight[22][39],
reservoir_weight[22][40],
reservoir_weight[22][41],
reservoir_weight[22][42],
reservoir_weight[22][43],
reservoir_weight[22][44],
reservoir_weight[22][45],
reservoir_weight[22][46],
reservoir_weight[22][47],
reservoir_weight[22][48],
reservoir_weight[22][49],
reservoir_weight[22][50],
reservoir_weight[22][51],
reservoir_weight[22][52],
reservoir_weight[22][53],
reservoir_weight[22][54],
reservoir_weight[22][55],
reservoir_weight[22][56],
reservoir_weight[22][57],
reservoir_weight[22][58],
reservoir_weight[22][59],
reservoir_weight[22][60],
reservoir_weight[22][61],
reservoir_weight[22][62],
reservoir_weight[22][63],
reservoir_weight[22][64],
reservoir_weight[22][65],
reservoir_weight[22][66],
reservoir_weight[22][67],
reservoir_weight[22][68],
reservoir_weight[22][69],
reservoir_weight[22][70],
reservoir_weight[22][71],
reservoir_weight[22][72],
reservoir_weight[22][73],
reservoir_weight[22][74],
reservoir_weight[22][75],
reservoir_weight[22][76],
reservoir_weight[22][77],
reservoir_weight[22][78],
reservoir_weight[22][79],
reservoir_weight[22][80],
reservoir_weight[22][81],
reservoir_weight[22][82],
reservoir_weight[22][83],
reservoir_weight[22][84],
reservoir_weight[22][85],
reservoir_weight[22][86],
reservoir_weight[22][87],
reservoir_weight[22][88],
reservoir_weight[22][89],
reservoir_weight[22][90],
reservoir_weight[22][91],
reservoir_weight[22][92],
reservoir_weight[22][93],
reservoir_weight[22][94],
reservoir_weight[22][95],
reservoir_weight[22][96],
reservoir_weight[22][97],
reservoir_weight[22][98],
reservoir_weight[22][99],
reservoir_weight[22][100],
reservoir_weight[22][101],
reservoir_weight[22][102],
reservoir_weight[22][103],
reservoir_weight[22][104],
reservoir_weight[22][105],
reservoir_weight[22][106],
reservoir_weight[22][107],
reservoir_weight[22][108],
reservoir_weight[22][109],
reservoir_weight[22][110],
reservoir_weight[22][111],
reservoir_weight[22][112],
reservoir_weight[22][113],
reservoir_weight[22][114],
reservoir_weight[22][115],
reservoir_weight[22][116],
reservoir_weight[22][117],
reservoir_weight[22][118],
reservoir_weight[22][119],
reservoir_weight[22][120],
reservoir_weight[22][121],
reservoir_weight[22][122],
reservoir_weight[22][123],
reservoir_weight[22][124],
reservoir_weight[22][125],
reservoir_weight[22][126],
reservoir_weight[22][127],
reservoir_weight[22][128],
reservoir_weight[22][129],
reservoir_weight[22][130],
reservoir_weight[22][131],
reservoir_weight[22][132],
reservoir_weight[22][133],
reservoir_weight[22][134],
reservoir_weight[22][135],
reservoir_weight[22][136],
reservoir_weight[22][137],
reservoir_weight[22][138],
reservoir_weight[22][139],
reservoir_weight[22][140],
reservoir_weight[22][141],
reservoir_weight[22][142],
reservoir_weight[22][143],
reservoir_weight[22][144],
reservoir_weight[22][145],
reservoir_weight[22][146],
reservoir_weight[22][147],
reservoir_weight[22][148],
reservoir_weight[22][149],
reservoir_weight[22][150],
reservoir_weight[22][151],
reservoir_weight[22][152],
reservoir_weight[22][153],
reservoir_weight[22][154],
reservoir_weight[22][155],
reservoir_weight[22][156],
reservoir_weight[22][157],
reservoir_weight[22][158],
reservoir_weight[22][159],
reservoir_weight[22][160],
reservoir_weight[22][161],
reservoir_weight[22][162],
reservoir_weight[22][163],
reservoir_weight[22][164],
reservoir_weight[22][165],
reservoir_weight[22][166],
reservoir_weight[22][167],
reservoir_weight[22][168],
reservoir_weight[22][169],
reservoir_weight[22][170],
reservoir_weight[22][171],
reservoir_weight[22][172],
reservoir_weight[22][173],
reservoir_weight[22][174],
reservoir_weight[22][175],
reservoir_weight[22][176],
reservoir_weight[22][177],
reservoir_weight[22][178],
reservoir_weight[22][179],
reservoir_weight[22][180],
reservoir_weight[22][181],
reservoir_weight[22][182],
reservoir_weight[22][183],
reservoir_weight[22][184],
reservoir_weight[22][185],
reservoir_weight[22][186],
reservoir_weight[22][187],
reservoir_weight[22][188],
reservoir_weight[22][189],
reservoir_weight[22][190],
reservoir_weight[22][191],
reservoir_weight[22][192],
reservoir_weight[22][193],
reservoir_weight[22][194],
reservoir_weight[22][195],
reservoir_weight[22][196],
reservoir_weight[22][197],
reservoir_weight[22][198],
reservoir_weight[22][199]
},
{reservoir_weight[23][0],
reservoir_weight[23][1],
reservoir_weight[23][2],
reservoir_weight[23][3],
reservoir_weight[23][4],
reservoir_weight[23][5],
reservoir_weight[23][6],
reservoir_weight[23][7],
reservoir_weight[23][8],
reservoir_weight[23][9],
reservoir_weight[23][10],
reservoir_weight[23][11],
reservoir_weight[23][12],
reservoir_weight[23][13],
reservoir_weight[23][14],
reservoir_weight[23][15],
reservoir_weight[23][16],
reservoir_weight[23][17],
reservoir_weight[23][18],
reservoir_weight[23][19],
reservoir_weight[23][20],
reservoir_weight[23][21],
reservoir_weight[23][22],
reservoir_weight[23][23],
reservoir_weight[23][24],
reservoir_weight[23][25],
reservoir_weight[23][26],
reservoir_weight[23][27],
reservoir_weight[23][28],
reservoir_weight[23][29],
reservoir_weight[23][30],
reservoir_weight[23][31],
reservoir_weight[23][32],
reservoir_weight[23][33],
reservoir_weight[23][34],
reservoir_weight[23][35],
reservoir_weight[23][36],
reservoir_weight[23][37],
reservoir_weight[23][38],
reservoir_weight[23][39],
reservoir_weight[23][40],
reservoir_weight[23][41],
reservoir_weight[23][42],
reservoir_weight[23][43],
reservoir_weight[23][44],
reservoir_weight[23][45],
reservoir_weight[23][46],
reservoir_weight[23][47],
reservoir_weight[23][48],
reservoir_weight[23][49],
reservoir_weight[23][50],
reservoir_weight[23][51],
reservoir_weight[23][52],
reservoir_weight[23][53],
reservoir_weight[23][54],
reservoir_weight[23][55],
reservoir_weight[23][56],
reservoir_weight[23][57],
reservoir_weight[23][58],
reservoir_weight[23][59],
reservoir_weight[23][60],
reservoir_weight[23][61],
reservoir_weight[23][62],
reservoir_weight[23][63],
reservoir_weight[23][64],
reservoir_weight[23][65],
reservoir_weight[23][66],
reservoir_weight[23][67],
reservoir_weight[23][68],
reservoir_weight[23][69],
reservoir_weight[23][70],
reservoir_weight[23][71],
reservoir_weight[23][72],
reservoir_weight[23][73],
reservoir_weight[23][74],
reservoir_weight[23][75],
reservoir_weight[23][76],
reservoir_weight[23][77],
reservoir_weight[23][78],
reservoir_weight[23][79],
reservoir_weight[23][80],
reservoir_weight[23][81],
reservoir_weight[23][82],
reservoir_weight[23][83],
reservoir_weight[23][84],
reservoir_weight[23][85],
reservoir_weight[23][86],
reservoir_weight[23][87],
reservoir_weight[23][88],
reservoir_weight[23][89],
reservoir_weight[23][90],
reservoir_weight[23][91],
reservoir_weight[23][92],
reservoir_weight[23][93],
reservoir_weight[23][94],
reservoir_weight[23][95],
reservoir_weight[23][96],
reservoir_weight[23][97],
reservoir_weight[23][98],
reservoir_weight[23][99],
reservoir_weight[23][100],
reservoir_weight[23][101],
reservoir_weight[23][102],
reservoir_weight[23][103],
reservoir_weight[23][104],
reservoir_weight[23][105],
reservoir_weight[23][106],
reservoir_weight[23][107],
reservoir_weight[23][108],
reservoir_weight[23][109],
reservoir_weight[23][110],
reservoir_weight[23][111],
reservoir_weight[23][112],
reservoir_weight[23][113],
reservoir_weight[23][114],
reservoir_weight[23][115],
reservoir_weight[23][116],
reservoir_weight[23][117],
reservoir_weight[23][118],
reservoir_weight[23][119],
reservoir_weight[23][120],
reservoir_weight[23][121],
reservoir_weight[23][122],
reservoir_weight[23][123],
reservoir_weight[23][124],
reservoir_weight[23][125],
reservoir_weight[23][126],
reservoir_weight[23][127],
reservoir_weight[23][128],
reservoir_weight[23][129],
reservoir_weight[23][130],
reservoir_weight[23][131],
reservoir_weight[23][132],
reservoir_weight[23][133],
reservoir_weight[23][134],
reservoir_weight[23][135],
reservoir_weight[23][136],
reservoir_weight[23][137],
reservoir_weight[23][138],
reservoir_weight[23][139],
reservoir_weight[23][140],
reservoir_weight[23][141],
reservoir_weight[23][142],
reservoir_weight[23][143],
reservoir_weight[23][144],
reservoir_weight[23][145],
reservoir_weight[23][146],
reservoir_weight[23][147],
reservoir_weight[23][148],
reservoir_weight[23][149],
reservoir_weight[23][150],
reservoir_weight[23][151],
reservoir_weight[23][152],
reservoir_weight[23][153],
reservoir_weight[23][154],
reservoir_weight[23][155],
reservoir_weight[23][156],
reservoir_weight[23][157],
reservoir_weight[23][158],
reservoir_weight[23][159],
reservoir_weight[23][160],
reservoir_weight[23][161],
reservoir_weight[23][162],
reservoir_weight[23][163],
reservoir_weight[23][164],
reservoir_weight[23][165],
reservoir_weight[23][166],
reservoir_weight[23][167],
reservoir_weight[23][168],
reservoir_weight[23][169],
reservoir_weight[23][170],
reservoir_weight[23][171],
reservoir_weight[23][172],
reservoir_weight[23][173],
reservoir_weight[23][174],
reservoir_weight[23][175],
reservoir_weight[23][176],
reservoir_weight[23][177],
reservoir_weight[23][178],
reservoir_weight[23][179],
reservoir_weight[23][180],
reservoir_weight[23][181],
reservoir_weight[23][182],
reservoir_weight[23][183],
reservoir_weight[23][184],
reservoir_weight[23][185],
reservoir_weight[23][186],
reservoir_weight[23][187],
reservoir_weight[23][188],
reservoir_weight[23][189],
reservoir_weight[23][190],
reservoir_weight[23][191],
reservoir_weight[23][192],
reservoir_weight[23][193],
reservoir_weight[23][194],
reservoir_weight[23][195],
reservoir_weight[23][196],
reservoir_weight[23][197],
reservoir_weight[23][198],
reservoir_weight[23][199]
},
{reservoir_weight[24][0],
reservoir_weight[24][1],
reservoir_weight[24][2],
reservoir_weight[24][3],
reservoir_weight[24][4],
reservoir_weight[24][5],
reservoir_weight[24][6],
reservoir_weight[24][7],
reservoir_weight[24][8],
reservoir_weight[24][9],
reservoir_weight[24][10],
reservoir_weight[24][11],
reservoir_weight[24][12],
reservoir_weight[24][13],
reservoir_weight[24][14],
reservoir_weight[24][15],
reservoir_weight[24][16],
reservoir_weight[24][17],
reservoir_weight[24][18],
reservoir_weight[24][19],
reservoir_weight[24][20],
reservoir_weight[24][21],
reservoir_weight[24][22],
reservoir_weight[24][23],
reservoir_weight[24][24],
reservoir_weight[24][25],
reservoir_weight[24][26],
reservoir_weight[24][27],
reservoir_weight[24][28],
reservoir_weight[24][29],
reservoir_weight[24][30],
reservoir_weight[24][31],
reservoir_weight[24][32],
reservoir_weight[24][33],
reservoir_weight[24][34],
reservoir_weight[24][35],
reservoir_weight[24][36],
reservoir_weight[24][37],
reservoir_weight[24][38],
reservoir_weight[24][39],
reservoir_weight[24][40],
reservoir_weight[24][41],
reservoir_weight[24][42],
reservoir_weight[24][43],
reservoir_weight[24][44],
reservoir_weight[24][45],
reservoir_weight[24][46],
reservoir_weight[24][47],
reservoir_weight[24][48],
reservoir_weight[24][49],
reservoir_weight[24][50],
reservoir_weight[24][51],
reservoir_weight[24][52],
reservoir_weight[24][53],
reservoir_weight[24][54],
reservoir_weight[24][55],
reservoir_weight[24][56],
reservoir_weight[24][57],
reservoir_weight[24][58],
reservoir_weight[24][59],
reservoir_weight[24][60],
reservoir_weight[24][61],
reservoir_weight[24][62],
reservoir_weight[24][63],
reservoir_weight[24][64],
reservoir_weight[24][65],
reservoir_weight[24][66],
reservoir_weight[24][67],
reservoir_weight[24][68],
reservoir_weight[24][69],
reservoir_weight[24][70],
reservoir_weight[24][71],
reservoir_weight[24][72],
reservoir_weight[24][73],
reservoir_weight[24][74],
reservoir_weight[24][75],
reservoir_weight[24][76],
reservoir_weight[24][77],
reservoir_weight[24][78],
reservoir_weight[24][79],
reservoir_weight[24][80],
reservoir_weight[24][81],
reservoir_weight[24][82],
reservoir_weight[24][83],
reservoir_weight[24][84],
reservoir_weight[24][85],
reservoir_weight[24][86],
reservoir_weight[24][87],
reservoir_weight[24][88],
reservoir_weight[24][89],
reservoir_weight[24][90],
reservoir_weight[24][91],
reservoir_weight[24][92],
reservoir_weight[24][93],
reservoir_weight[24][94],
reservoir_weight[24][95],
reservoir_weight[24][96],
reservoir_weight[24][97],
reservoir_weight[24][98],
reservoir_weight[24][99],
reservoir_weight[24][100],
reservoir_weight[24][101],
reservoir_weight[24][102],
reservoir_weight[24][103],
reservoir_weight[24][104],
reservoir_weight[24][105],
reservoir_weight[24][106],
reservoir_weight[24][107],
reservoir_weight[24][108],
reservoir_weight[24][109],
reservoir_weight[24][110],
reservoir_weight[24][111],
reservoir_weight[24][112],
reservoir_weight[24][113],
reservoir_weight[24][114],
reservoir_weight[24][115],
reservoir_weight[24][116],
reservoir_weight[24][117],
reservoir_weight[24][118],
reservoir_weight[24][119],
reservoir_weight[24][120],
reservoir_weight[24][121],
reservoir_weight[24][122],
reservoir_weight[24][123],
reservoir_weight[24][124],
reservoir_weight[24][125],
reservoir_weight[24][126],
reservoir_weight[24][127],
reservoir_weight[24][128],
reservoir_weight[24][129],
reservoir_weight[24][130],
reservoir_weight[24][131],
reservoir_weight[24][132],
reservoir_weight[24][133],
reservoir_weight[24][134],
reservoir_weight[24][135],
reservoir_weight[24][136],
reservoir_weight[24][137],
reservoir_weight[24][138],
reservoir_weight[24][139],
reservoir_weight[24][140],
reservoir_weight[24][141],
reservoir_weight[24][142],
reservoir_weight[24][143],
reservoir_weight[24][144],
reservoir_weight[24][145],
reservoir_weight[24][146],
reservoir_weight[24][147],
reservoir_weight[24][148],
reservoir_weight[24][149],
reservoir_weight[24][150],
reservoir_weight[24][151],
reservoir_weight[24][152],
reservoir_weight[24][153],
reservoir_weight[24][154],
reservoir_weight[24][155],
reservoir_weight[24][156],
reservoir_weight[24][157],
reservoir_weight[24][158],
reservoir_weight[24][159],
reservoir_weight[24][160],
reservoir_weight[24][161],
reservoir_weight[24][162],
reservoir_weight[24][163],
reservoir_weight[24][164],
reservoir_weight[24][165],
reservoir_weight[24][166],
reservoir_weight[24][167],
reservoir_weight[24][168],
reservoir_weight[24][169],
reservoir_weight[24][170],
reservoir_weight[24][171],
reservoir_weight[24][172],
reservoir_weight[24][173],
reservoir_weight[24][174],
reservoir_weight[24][175],
reservoir_weight[24][176],
reservoir_weight[24][177],
reservoir_weight[24][178],
reservoir_weight[24][179],
reservoir_weight[24][180],
reservoir_weight[24][181],
reservoir_weight[24][182],
reservoir_weight[24][183],
reservoir_weight[24][184],
reservoir_weight[24][185],
reservoir_weight[24][186],
reservoir_weight[24][187],
reservoir_weight[24][188],
reservoir_weight[24][189],
reservoir_weight[24][190],
reservoir_weight[24][191],
reservoir_weight[24][192],
reservoir_weight[24][193],
reservoir_weight[24][194],
reservoir_weight[24][195],
reservoir_weight[24][196],
reservoir_weight[24][197],
reservoir_weight[24][198],
reservoir_weight[24][199]
},
{reservoir_weight[25][0],
reservoir_weight[25][1],
reservoir_weight[25][2],
reservoir_weight[25][3],
reservoir_weight[25][4],
reservoir_weight[25][5],
reservoir_weight[25][6],
reservoir_weight[25][7],
reservoir_weight[25][8],
reservoir_weight[25][9],
reservoir_weight[25][10],
reservoir_weight[25][11],
reservoir_weight[25][12],
reservoir_weight[25][13],
reservoir_weight[25][14],
reservoir_weight[25][15],
reservoir_weight[25][16],
reservoir_weight[25][17],
reservoir_weight[25][18],
reservoir_weight[25][19],
reservoir_weight[25][20],
reservoir_weight[25][21],
reservoir_weight[25][22],
reservoir_weight[25][23],
reservoir_weight[25][24],
reservoir_weight[25][25],
reservoir_weight[25][26],
reservoir_weight[25][27],
reservoir_weight[25][28],
reservoir_weight[25][29],
reservoir_weight[25][30],
reservoir_weight[25][31],
reservoir_weight[25][32],
reservoir_weight[25][33],
reservoir_weight[25][34],
reservoir_weight[25][35],
reservoir_weight[25][36],
reservoir_weight[25][37],
reservoir_weight[25][38],
reservoir_weight[25][39],
reservoir_weight[25][40],
reservoir_weight[25][41],
reservoir_weight[25][42],
reservoir_weight[25][43],
reservoir_weight[25][44],
reservoir_weight[25][45],
reservoir_weight[25][46],
reservoir_weight[25][47],
reservoir_weight[25][48],
reservoir_weight[25][49],
reservoir_weight[25][50],
reservoir_weight[25][51],
reservoir_weight[25][52],
reservoir_weight[25][53],
reservoir_weight[25][54],
reservoir_weight[25][55],
reservoir_weight[25][56],
reservoir_weight[25][57],
reservoir_weight[25][58],
reservoir_weight[25][59],
reservoir_weight[25][60],
reservoir_weight[25][61],
reservoir_weight[25][62],
reservoir_weight[25][63],
reservoir_weight[25][64],
reservoir_weight[25][65],
reservoir_weight[25][66],
reservoir_weight[25][67],
reservoir_weight[25][68],
reservoir_weight[25][69],
reservoir_weight[25][70],
reservoir_weight[25][71],
reservoir_weight[25][72],
reservoir_weight[25][73],
reservoir_weight[25][74],
reservoir_weight[25][75],
reservoir_weight[25][76],
reservoir_weight[25][77],
reservoir_weight[25][78],
reservoir_weight[25][79],
reservoir_weight[25][80],
reservoir_weight[25][81],
reservoir_weight[25][82],
reservoir_weight[25][83],
reservoir_weight[25][84],
reservoir_weight[25][85],
reservoir_weight[25][86],
reservoir_weight[25][87],
reservoir_weight[25][88],
reservoir_weight[25][89],
reservoir_weight[25][90],
reservoir_weight[25][91],
reservoir_weight[25][92],
reservoir_weight[25][93],
reservoir_weight[25][94],
reservoir_weight[25][95],
reservoir_weight[25][96],
reservoir_weight[25][97],
reservoir_weight[25][98],
reservoir_weight[25][99],
reservoir_weight[25][100],
reservoir_weight[25][101],
reservoir_weight[25][102],
reservoir_weight[25][103],
reservoir_weight[25][104],
reservoir_weight[25][105],
reservoir_weight[25][106],
reservoir_weight[25][107],
reservoir_weight[25][108],
reservoir_weight[25][109],
reservoir_weight[25][110],
reservoir_weight[25][111],
reservoir_weight[25][112],
reservoir_weight[25][113],
reservoir_weight[25][114],
reservoir_weight[25][115],
reservoir_weight[25][116],
reservoir_weight[25][117],
reservoir_weight[25][118],
reservoir_weight[25][119],
reservoir_weight[25][120],
reservoir_weight[25][121],
reservoir_weight[25][122],
reservoir_weight[25][123],
reservoir_weight[25][124],
reservoir_weight[25][125],
reservoir_weight[25][126],
reservoir_weight[25][127],
reservoir_weight[25][128],
reservoir_weight[25][129],
reservoir_weight[25][130],
reservoir_weight[25][131],
reservoir_weight[25][132],
reservoir_weight[25][133],
reservoir_weight[25][134],
reservoir_weight[25][135],
reservoir_weight[25][136],
reservoir_weight[25][137],
reservoir_weight[25][138],
reservoir_weight[25][139],
reservoir_weight[25][140],
reservoir_weight[25][141],
reservoir_weight[25][142],
reservoir_weight[25][143],
reservoir_weight[25][144],
reservoir_weight[25][145],
reservoir_weight[25][146],
reservoir_weight[25][147],
reservoir_weight[25][148],
reservoir_weight[25][149],
reservoir_weight[25][150],
reservoir_weight[25][151],
reservoir_weight[25][152],
reservoir_weight[25][153],
reservoir_weight[25][154],
reservoir_weight[25][155],
reservoir_weight[25][156],
reservoir_weight[25][157],
reservoir_weight[25][158],
reservoir_weight[25][159],
reservoir_weight[25][160],
reservoir_weight[25][161],
reservoir_weight[25][162],
reservoir_weight[25][163],
reservoir_weight[25][164],
reservoir_weight[25][165],
reservoir_weight[25][166],
reservoir_weight[25][167],
reservoir_weight[25][168],
reservoir_weight[25][169],
reservoir_weight[25][170],
reservoir_weight[25][171],
reservoir_weight[25][172],
reservoir_weight[25][173],
reservoir_weight[25][174],
reservoir_weight[25][175],
reservoir_weight[25][176],
reservoir_weight[25][177],
reservoir_weight[25][178],
reservoir_weight[25][179],
reservoir_weight[25][180],
reservoir_weight[25][181],
reservoir_weight[25][182],
reservoir_weight[25][183],
reservoir_weight[25][184],
reservoir_weight[25][185],
reservoir_weight[25][186],
reservoir_weight[25][187],
reservoir_weight[25][188],
reservoir_weight[25][189],
reservoir_weight[25][190],
reservoir_weight[25][191],
reservoir_weight[25][192],
reservoir_weight[25][193],
reservoir_weight[25][194],
reservoir_weight[25][195],
reservoir_weight[25][196],
reservoir_weight[25][197],
reservoir_weight[25][198],
reservoir_weight[25][199]
},
{reservoir_weight[26][0],
reservoir_weight[26][1],
reservoir_weight[26][2],
reservoir_weight[26][3],
reservoir_weight[26][4],
reservoir_weight[26][5],
reservoir_weight[26][6],
reservoir_weight[26][7],
reservoir_weight[26][8],
reservoir_weight[26][9],
reservoir_weight[26][10],
reservoir_weight[26][11],
reservoir_weight[26][12],
reservoir_weight[26][13],
reservoir_weight[26][14],
reservoir_weight[26][15],
reservoir_weight[26][16],
reservoir_weight[26][17],
reservoir_weight[26][18],
reservoir_weight[26][19],
reservoir_weight[26][20],
reservoir_weight[26][21],
reservoir_weight[26][22],
reservoir_weight[26][23],
reservoir_weight[26][24],
reservoir_weight[26][25],
reservoir_weight[26][26],
reservoir_weight[26][27],
reservoir_weight[26][28],
reservoir_weight[26][29],
reservoir_weight[26][30],
reservoir_weight[26][31],
reservoir_weight[26][32],
reservoir_weight[26][33],
reservoir_weight[26][34],
reservoir_weight[26][35],
reservoir_weight[26][36],
reservoir_weight[26][37],
reservoir_weight[26][38],
reservoir_weight[26][39],
reservoir_weight[26][40],
reservoir_weight[26][41],
reservoir_weight[26][42],
reservoir_weight[26][43],
reservoir_weight[26][44],
reservoir_weight[26][45],
reservoir_weight[26][46],
reservoir_weight[26][47],
reservoir_weight[26][48],
reservoir_weight[26][49],
reservoir_weight[26][50],
reservoir_weight[26][51],
reservoir_weight[26][52],
reservoir_weight[26][53],
reservoir_weight[26][54],
reservoir_weight[26][55],
reservoir_weight[26][56],
reservoir_weight[26][57],
reservoir_weight[26][58],
reservoir_weight[26][59],
reservoir_weight[26][60],
reservoir_weight[26][61],
reservoir_weight[26][62],
reservoir_weight[26][63],
reservoir_weight[26][64],
reservoir_weight[26][65],
reservoir_weight[26][66],
reservoir_weight[26][67],
reservoir_weight[26][68],
reservoir_weight[26][69],
reservoir_weight[26][70],
reservoir_weight[26][71],
reservoir_weight[26][72],
reservoir_weight[26][73],
reservoir_weight[26][74],
reservoir_weight[26][75],
reservoir_weight[26][76],
reservoir_weight[26][77],
reservoir_weight[26][78],
reservoir_weight[26][79],
reservoir_weight[26][80],
reservoir_weight[26][81],
reservoir_weight[26][82],
reservoir_weight[26][83],
reservoir_weight[26][84],
reservoir_weight[26][85],
reservoir_weight[26][86],
reservoir_weight[26][87],
reservoir_weight[26][88],
reservoir_weight[26][89],
reservoir_weight[26][90],
reservoir_weight[26][91],
reservoir_weight[26][92],
reservoir_weight[26][93],
reservoir_weight[26][94],
reservoir_weight[26][95],
reservoir_weight[26][96],
reservoir_weight[26][97],
reservoir_weight[26][98],
reservoir_weight[26][99],
reservoir_weight[26][100],
reservoir_weight[26][101],
reservoir_weight[26][102],
reservoir_weight[26][103],
reservoir_weight[26][104],
reservoir_weight[26][105],
reservoir_weight[26][106],
reservoir_weight[26][107],
reservoir_weight[26][108],
reservoir_weight[26][109],
reservoir_weight[26][110],
reservoir_weight[26][111],
reservoir_weight[26][112],
reservoir_weight[26][113],
reservoir_weight[26][114],
reservoir_weight[26][115],
reservoir_weight[26][116],
reservoir_weight[26][117],
reservoir_weight[26][118],
reservoir_weight[26][119],
reservoir_weight[26][120],
reservoir_weight[26][121],
reservoir_weight[26][122],
reservoir_weight[26][123],
reservoir_weight[26][124],
reservoir_weight[26][125],
reservoir_weight[26][126],
reservoir_weight[26][127],
reservoir_weight[26][128],
reservoir_weight[26][129],
reservoir_weight[26][130],
reservoir_weight[26][131],
reservoir_weight[26][132],
reservoir_weight[26][133],
reservoir_weight[26][134],
reservoir_weight[26][135],
reservoir_weight[26][136],
reservoir_weight[26][137],
reservoir_weight[26][138],
reservoir_weight[26][139],
reservoir_weight[26][140],
reservoir_weight[26][141],
reservoir_weight[26][142],
reservoir_weight[26][143],
reservoir_weight[26][144],
reservoir_weight[26][145],
reservoir_weight[26][146],
reservoir_weight[26][147],
reservoir_weight[26][148],
reservoir_weight[26][149],
reservoir_weight[26][150],
reservoir_weight[26][151],
reservoir_weight[26][152],
reservoir_weight[26][153],
reservoir_weight[26][154],
reservoir_weight[26][155],
reservoir_weight[26][156],
reservoir_weight[26][157],
reservoir_weight[26][158],
reservoir_weight[26][159],
reservoir_weight[26][160],
reservoir_weight[26][161],
reservoir_weight[26][162],
reservoir_weight[26][163],
reservoir_weight[26][164],
reservoir_weight[26][165],
reservoir_weight[26][166],
reservoir_weight[26][167],
reservoir_weight[26][168],
reservoir_weight[26][169],
reservoir_weight[26][170],
reservoir_weight[26][171],
reservoir_weight[26][172],
reservoir_weight[26][173],
reservoir_weight[26][174],
reservoir_weight[26][175],
reservoir_weight[26][176],
reservoir_weight[26][177],
reservoir_weight[26][178],
reservoir_weight[26][179],
reservoir_weight[26][180],
reservoir_weight[26][181],
reservoir_weight[26][182],
reservoir_weight[26][183],
reservoir_weight[26][184],
reservoir_weight[26][185],
reservoir_weight[26][186],
reservoir_weight[26][187],
reservoir_weight[26][188],
reservoir_weight[26][189],
reservoir_weight[26][190],
reservoir_weight[26][191],
reservoir_weight[26][192],
reservoir_weight[26][193],
reservoir_weight[26][194],
reservoir_weight[26][195],
reservoir_weight[26][196],
reservoir_weight[26][197],
reservoir_weight[26][198],
reservoir_weight[26][199]
},
{reservoir_weight[27][0],
reservoir_weight[27][1],
reservoir_weight[27][2],
reservoir_weight[27][3],
reservoir_weight[27][4],
reservoir_weight[27][5],
reservoir_weight[27][6],
reservoir_weight[27][7],
reservoir_weight[27][8],
reservoir_weight[27][9],
reservoir_weight[27][10],
reservoir_weight[27][11],
reservoir_weight[27][12],
reservoir_weight[27][13],
reservoir_weight[27][14],
reservoir_weight[27][15],
reservoir_weight[27][16],
reservoir_weight[27][17],
reservoir_weight[27][18],
reservoir_weight[27][19],
reservoir_weight[27][20],
reservoir_weight[27][21],
reservoir_weight[27][22],
reservoir_weight[27][23],
reservoir_weight[27][24],
reservoir_weight[27][25],
reservoir_weight[27][26],
reservoir_weight[27][27],
reservoir_weight[27][28],
reservoir_weight[27][29],
reservoir_weight[27][30],
reservoir_weight[27][31],
reservoir_weight[27][32],
reservoir_weight[27][33],
reservoir_weight[27][34],
reservoir_weight[27][35],
reservoir_weight[27][36],
reservoir_weight[27][37],
reservoir_weight[27][38],
reservoir_weight[27][39],
reservoir_weight[27][40],
reservoir_weight[27][41],
reservoir_weight[27][42],
reservoir_weight[27][43],
reservoir_weight[27][44],
reservoir_weight[27][45],
reservoir_weight[27][46],
reservoir_weight[27][47],
reservoir_weight[27][48],
reservoir_weight[27][49],
reservoir_weight[27][50],
reservoir_weight[27][51],
reservoir_weight[27][52],
reservoir_weight[27][53],
reservoir_weight[27][54],
reservoir_weight[27][55],
reservoir_weight[27][56],
reservoir_weight[27][57],
reservoir_weight[27][58],
reservoir_weight[27][59],
reservoir_weight[27][60],
reservoir_weight[27][61],
reservoir_weight[27][62],
reservoir_weight[27][63],
reservoir_weight[27][64],
reservoir_weight[27][65],
reservoir_weight[27][66],
reservoir_weight[27][67],
reservoir_weight[27][68],
reservoir_weight[27][69],
reservoir_weight[27][70],
reservoir_weight[27][71],
reservoir_weight[27][72],
reservoir_weight[27][73],
reservoir_weight[27][74],
reservoir_weight[27][75],
reservoir_weight[27][76],
reservoir_weight[27][77],
reservoir_weight[27][78],
reservoir_weight[27][79],
reservoir_weight[27][80],
reservoir_weight[27][81],
reservoir_weight[27][82],
reservoir_weight[27][83],
reservoir_weight[27][84],
reservoir_weight[27][85],
reservoir_weight[27][86],
reservoir_weight[27][87],
reservoir_weight[27][88],
reservoir_weight[27][89],
reservoir_weight[27][90],
reservoir_weight[27][91],
reservoir_weight[27][92],
reservoir_weight[27][93],
reservoir_weight[27][94],
reservoir_weight[27][95],
reservoir_weight[27][96],
reservoir_weight[27][97],
reservoir_weight[27][98],
reservoir_weight[27][99],
reservoir_weight[27][100],
reservoir_weight[27][101],
reservoir_weight[27][102],
reservoir_weight[27][103],
reservoir_weight[27][104],
reservoir_weight[27][105],
reservoir_weight[27][106],
reservoir_weight[27][107],
reservoir_weight[27][108],
reservoir_weight[27][109],
reservoir_weight[27][110],
reservoir_weight[27][111],
reservoir_weight[27][112],
reservoir_weight[27][113],
reservoir_weight[27][114],
reservoir_weight[27][115],
reservoir_weight[27][116],
reservoir_weight[27][117],
reservoir_weight[27][118],
reservoir_weight[27][119],
reservoir_weight[27][120],
reservoir_weight[27][121],
reservoir_weight[27][122],
reservoir_weight[27][123],
reservoir_weight[27][124],
reservoir_weight[27][125],
reservoir_weight[27][126],
reservoir_weight[27][127],
reservoir_weight[27][128],
reservoir_weight[27][129],
reservoir_weight[27][130],
reservoir_weight[27][131],
reservoir_weight[27][132],
reservoir_weight[27][133],
reservoir_weight[27][134],
reservoir_weight[27][135],
reservoir_weight[27][136],
reservoir_weight[27][137],
reservoir_weight[27][138],
reservoir_weight[27][139],
reservoir_weight[27][140],
reservoir_weight[27][141],
reservoir_weight[27][142],
reservoir_weight[27][143],
reservoir_weight[27][144],
reservoir_weight[27][145],
reservoir_weight[27][146],
reservoir_weight[27][147],
reservoir_weight[27][148],
reservoir_weight[27][149],
reservoir_weight[27][150],
reservoir_weight[27][151],
reservoir_weight[27][152],
reservoir_weight[27][153],
reservoir_weight[27][154],
reservoir_weight[27][155],
reservoir_weight[27][156],
reservoir_weight[27][157],
reservoir_weight[27][158],
reservoir_weight[27][159],
reservoir_weight[27][160],
reservoir_weight[27][161],
reservoir_weight[27][162],
reservoir_weight[27][163],
reservoir_weight[27][164],
reservoir_weight[27][165],
reservoir_weight[27][166],
reservoir_weight[27][167],
reservoir_weight[27][168],
reservoir_weight[27][169],
reservoir_weight[27][170],
reservoir_weight[27][171],
reservoir_weight[27][172],
reservoir_weight[27][173],
reservoir_weight[27][174],
reservoir_weight[27][175],
reservoir_weight[27][176],
reservoir_weight[27][177],
reservoir_weight[27][178],
reservoir_weight[27][179],
reservoir_weight[27][180],
reservoir_weight[27][181],
reservoir_weight[27][182],
reservoir_weight[27][183],
reservoir_weight[27][184],
reservoir_weight[27][185],
reservoir_weight[27][186],
reservoir_weight[27][187],
reservoir_weight[27][188],
reservoir_weight[27][189],
reservoir_weight[27][190],
reservoir_weight[27][191],
reservoir_weight[27][192],
reservoir_weight[27][193],
reservoir_weight[27][194],
reservoir_weight[27][195],
reservoir_weight[27][196],
reservoir_weight[27][197],
reservoir_weight[27][198],
reservoir_weight[27][199]
},
{reservoir_weight[28][0],
reservoir_weight[28][1],
reservoir_weight[28][2],
reservoir_weight[28][3],
reservoir_weight[28][4],
reservoir_weight[28][5],
reservoir_weight[28][6],
reservoir_weight[28][7],
reservoir_weight[28][8],
reservoir_weight[28][9],
reservoir_weight[28][10],
reservoir_weight[28][11],
reservoir_weight[28][12],
reservoir_weight[28][13],
reservoir_weight[28][14],
reservoir_weight[28][15],
reservoir_weight[28][16],
reservoir_weight[28][17],
reservoir_weight[28][18],
reservoir_weight[28][19],
reservoir_weight[28][20],
reservoir_weight[28][21],
reservoir_weight[28][22],
reservoir_weight[28][23],
reservoir_weight[28][24],
reservoir_weight[28][25],
reservoir_weight[28][26],
reservoir_weight[28][27],
reservoir_weight[28][28],
reservoir_weight[28][29],
reservoir_weight[28][30],
reservoir_weight[28][31],
reservoir_weight[28][32],
reservoir_weight[28][33],
reservoir_weight[28][34],
reservoir_weight[28][35],
reservoir_weight[28][36],
reservoir_weight[28][37],
reservoir_weight[28][38],
reservoir_weight[28][39],
reservoir_weight[28][40],
reservoir_weight[28][41],
reservoir_weight[28][42],
reservoir_weight[28][43],
reservoir_weight[28][44],
reservoir_weight[28][45],
reservoir_weight[28][46],
reservoir_weight[28][47],
reservoir_weight[28][48],
reservoir_weight[28][49],
reservoir_weight[28][50],
reservoir_weight[28][51],
reservoir_weight[28][52],
reservoir_weight[28][53],
reservoir_weight[28][54],
reservoir_weight[28][55],
reservoir_weight[28][56],
reservoir_weight[28][57],
reservoir_weight[28][58],
reservoir_weight[28][59],
reservoir_weight[28][60],
reservoir_weight[28][61],
reservoir_weight[28][62],
reservoir_weight[28][63],
reservoir_weight[28][64],
reservoir_weight[28][65],
reservoir_weight[28][66],
reservoir_weight[28][67],
reservoir_weight[28][68],
reservoir_weight[28][69],
reservoir_weight[28][70],
reservoir_weight[28][71],
reservoir_weight[28][72],
reservoir_weight[28][73],
reservoir_weight[28][74],
reservoir_weight[28][75],
reservoir_weight[28][76],
reservoir_weight[28][77],
reservoir_weight[28][78],
reservoir_weight[28][79],
reservoir_weight[28][80],
reservoir_weight[28][81],
reservoir_weight[28][82],
reservoir_weight[28][83],
reservoir_weight[28][84],
reservoir_weight[28][85],
reservoir_weight[28][86],
reservoir_weight[28][87],
reservoir_weight[28][88],
reservoir_weight[28][89],
reservoir_weight[28][90],
reservoir_weight[28][91],
reservoir_weight[28][92],
reservoir_weight[28][93],
reservoir_weight[28][94],
reservoir_weight[28][95],
reservoir_weight[28][96],
reservoir_weight[28][97],
reservoir_weight[28][98],
reservoir_weight[28][99],
reservoir_weight[28][100],
reservoir_weight[28][101],
reservoir_weight[28][102],
reservoir_weight[28][103],
reservoir_weight[28][104],
reservoir_weight[28][105],
reservoir_weight[28][106],
reservoir_weight[28][107],
reservoir_weight[28][108],
reservoir_weight[28][109],
reservoir_weight[28][110],
reservoir_weight[28][111],
reservoir_weight[28][112],
reservoir_weight[28][113],
reservoir_weight[28][114],
reservoir_weight[28][115],
reservoir_weight[28][116],
reservoir_weight[28][117],
reservoir_weight[28][118],
reservoir_weight[28][119],
reservoir_weight[28][120],
reservoir_weight[28][121],
reservoir_weight[28][122],
reservoir_weight[28][123],
reservoir_weight[28][124],
reservoir_weight[28][125],
reservoir_weight[28][126],
reservoir_weight[28][127],
reservoir_weight[28][128],
reservoir_weight[28][129],
reservoir_weight[28][130],
reservoir_weight[28][131],
reservoir_weight[28][132],
reservoir_weight[28][133],
reservoir_weight[28][134],
reservoir_weight[28][135],
reservoir_weight[28][136],
reservoir_weight[28][137],
reservoir_weight[28][138],
reservoir_weight[28][139],
reservoir_weight[28][140],
reservoir_weight[28][141],
reservoir_weight[28][142],
reservoir_weight[28][143],
reservoir_weight[28][144],
reservoir_weight[28][145],
reservoir_weight[28][146],
reservoir_weight[28][147],
reservoir_weight[28][148],
reservoir_weight[28][149],
reservoir_weight[28][150],
reservoir_weight[28][151],
reservoir_weight[28][152],
reservoir_weight[28][153],
reservoir_weight[28][154],
reservoir_weight[28][155],
reservoir_weight[28][156],
reservoir_weight[28][157],
reservoir_weight[28][158],
reservoir_weight[28][159],
reservoir_weight[28][160],
reservoir_weight[28][161],
reservoir_weight[28][162],
reservoir_weight[28][163],
reservoir_weight[28][164],
reservoir_weight[28][165],
reservoir_weight[28][166],
reservoir_weight[28][167],
reservoir_weight[28][168],
reservoir_weight[28][169],
reservoir_weight[28][170],
reservoir_weight[28][171],
reservoir_weight[28][172],
reservoir_weight[28][173],
reservoir_weight[28][174],
reservoir_weight[28][175],
reservoir_weight[28][176],
reservoir_weight[28][177],
reservoir_weight[28][178],
reservoir_weight[28][179],
reservoir_weight[28][180],
reservoir_weight[28][181],
reservoir_weight[28][182],
reservoir_weight[28][183],
reservoir_weight[28][184],
reservoir_weight[28][185],
reservoir_weight[28][186],
reservoir_weight[28][187],
reservoir_weight[28][188],
reservoir_weight[28][189],
reservoir_weight[28][190],
reservoir_weight[28][191],
reservoir_weight[28][192],
reservoir_weight[28][193],
reservoir_weight[28][194],
reservoir_weight[28][195],
reservoir_weight[28][196],
reservoir_weight[28][197],
reservoir_weight[28][198],
reservoir_weight[28][199]
},
{reservoir_weight[29][0],
reservoir_weight[29][1],
reservoir_weight[29][2],
reservoir_weight[29][3],
reservoir_weight[29][4],
reservoir_weight[29][5],
reservoir_weight[29][6],
reservoir_weight[29][7],
reservoir_weight[29][8],
reservoir_weight[29][9],
reservoir_weight[29][10],
reservoir_weight[29][11],
reservoir_weight[29][12],
reservoir_weight[29][13],
reservoir_weight[29][14],
reservoir_weight[29][15],
reservoir_weight[29][16],
reservoir_weight[29][17],
reservoir_weight[29][18],
reservoir_weight[29][19],
reservoir_weight[29][20],
reservoir_weight[29][21],
reservoir_weight[29][22],
reservoir_weight[29][23],
reservoir_weight[29][24],
reservoir_weight[29][25],
reservoir_weight[29][26],
reservoir_weight[29][27],
reservoir_weight[29][28],
reservoir_weight[29][29],
reservoir_weight[29][30],
reservoir_weight[29][31],
reservoir_weight[29][32],
reservoir_weight[29][33],
reservoir_weight[29][34],
reservoir_weight[29][35],
reservoir_weight[29][36],
reservoir_weight[29][37],
reservoir_weight[29][38],
reservoir_weight[29][39],
reservoir_weight[29][40],
reservoir_weight[29][41],
reservoir_weight[29][42],
reservoir_weight[29][43],
reservoir_weight[29][44],
reservoir_weight[29][45],
reservoir_weight[29][46],
reservoir_weight[29][47],
reservoir_weight[29][48],
reservoir_weight[29][49],
reservoir_weight[29][50],
reservoir_weight[29][51],
reservoir_weight[29][52],
reservoir_weight[29][53],
reservoir_weight[29][54],
reservoir_weight[29][55],
reservoir_weight[29][56],
reservoir_weight[29][57],
reservoir_weight[29][58],
reservoir_weight[29][59],
reservoir_weight[29][60],
reservoir_weight[29][61],
reservoir_weight[29][62],
reservoir_weight[29][63],
reservoir_weight[29][64],
reservoir_weight[29][65],
reservoir_weight[29][66],
reservoir_weight[29][67],
reservoir_weight[29][68],
reservoir_weight[29][69],
reservoir_weight[29][70],
reservoir_weight[29][71],
reservoir_weight[29][72],
reservoir_weight[29][73],
reservoir_weight[29][74],
reservoir_weight[29][75],
reservoir_weight[29][76],
reservoir_weight[29][77],
reservoir_weight[29][78],
reservoir_weight[29][79],
reservoir_weight[29][80],
reservoir_weight[29][81],
reservoir_weight[29][82],
reservoir_weight[29][83],
reservoir_weight[29][84],
reservoir_weight[29][85],
reservoir_weight[29][86],
reservoir_weight[29][87],
reservoir_weight[29][88],
reservoir_weight[29][89],
reservoir_weight[29][90],
reservoir_weight[29][91],
reservoir_weight[29][92],
reservoir_weight[29][93],
reservoir_weight[29][94],
reservoir_weight[29][95],
reservoir_weight[29][96],
reservoir_weight[29][97],
reservoir_weight[29][98],
reservoir_weight[29][99],
reservoir_weight[29][100],
reservoir_weight[29][101],
reservoir_weight[29][102],
reservoir_weight[29][103],
reservoir_weight[29][104],
reservoir_weight[29][105],
reservoir_weight[29][106],
reservoir_weight[29][107],
reservoir_weight[29][108],
reservoir_weight[29][109],
reservoir_weight[29][110],
reservoir_weight[29][111],
reservoir_weight[29][112],
reservoir_weight[29][113],
reservoir_weight[29][114],
reservoir_weight[29][115],
reservoir_weight[29][116],
reservoir_weight[29][117],
reservoir_weight[29][118],
reservoir_weight[29][119],
reservoir_weight[29][120],
reservoir_weight[29][121],
reservoir_weight[29][122],
reservoir_weight[29][123],
reservoir_weight[29][124],
reservoir_weight[29][125],
reservoir_weight[29][126],
reservoir_weight[29][127],
reservoir_weight[29][128],
reservoir_weight[29][129],
reservoir_weight[29][130],
reservoir_weight[29][131],
reservoir_weight[29][132],
reservoir_weight[29][133],
reservoir_weight[29][134],
reservoir_weight[29][135],
reservoir_weight[29][136],
reservoir_weight[29][137],
reservoir_weight[29][138],
reservoir_weight[29][139],
reservoir_weight[29][140],
reservoir_weight[29][141],
reservoir_weight[29][142],
reservoir_weight[29][143],
reservoir_weight[29][144],
reservoir_weight[29][145],
reservoir_weight[29][146],
reservoir_weight[29][147],
reservoir_weight[29][148],
reservoir_weight[29][149],
reservoir_weight[29][150],
reservoir_weight[29][151],
reservoir_weight[29][152],
reservoir_weight[29][153],
reservoir_weight[29][154],
reservoir_weight[29][155],
reservoir_weight[29][156],
reservoir_weight[29][157],
reservoir_weight[29][158],
reservoir_weight[29][159],
reservoir_weight[29][160],
reservoir_weight[29][161],
reservoir_weight[29][162],
reservoir_weight[29][163],
reservoir_weight[29][164],
reservoir_weight[29][165],
reservoir_weight[29][166],
reservoir_weight[29][167],
reservoir_weight[29][168],
reservoir_weight[29][169],
reservoir_weight[29][170],
reservoir_weight[29][171],
reservoir_weight[29][172],
reservoir_weight[29][173],
reservoir_weight[29][174],
reservoir_weight[29][175],
reservoir_weight[29][176],
reservoir_weight[29][177],
reservoir_weight[29][178],
reservoir_weight[29][179],
reservoir_weight[29][180],
reservoir_weight[29][181],
reservoir_weight[29][182],
reservoir_weight[29][183],
reservoir_weight[29][184],
reservoir_weight[29][185],
reservoir_weight[29][186],
reservoir_weight[29][187],
reservoir_weight[29][188],
reservoir_weight[29][189],
reservoir_weight[29][190],
reservoir_weight[29][191],
reservoir_weight[29][192],
reservoir_weight[29][193],
reservoir_weight[29][194],
reservoir_weight[29][195],
reservoir_weight[29][196],
reservoir_weight[29][197],
reservoir_weight[29][198],
reservoir_weight[29][199]
},
{reservoir_weight[30][0],
reservoir_weight[30][1],
reservoir_weight[30][2],
reservoir_weight[30][3],
reservoir_weight[30][4],
reservoir_weight[30][5],
reservoir_weight[30][6],
reservoir_weight[30][7],
reservoir_weight[30][8],
reservoir_weight[30][9],
reservoir_weight[30][10],
reservoir_weight[30][11],
reservoir_weight[30][12],
reservoir_weight[30][13],
reservoir_weight[30][14],
reservoir_weight[30][15],
reservoir_weight[30][16],
reservoir_weight[30][17],
reservoir_weight[30][18],
reservoir_weight[30][19],
reservoir_weight[30][20],
reservoir_weight[30][21],
reservoir_weight[30][22],
reservoir_weight[30][23],
reservoir_weight[30][24],
reservoir_weight[30][25],
reservoir_weight[30][26],
reservoir_weight[30][27],
reservoir_weight[30][28],
reservoir_weight[30][29],
reservoir_weight[30][30],
reservoir_weight[30][31],
reservoir_weight[30][32],
reservoir_weight[30][33],
reservoir_weight[30][34],
reservoir_weight[30][35],
reservoir_weight[30][36],
reservoir_weight[30][37],
reservoir_weight[30][38],
reservoir_weight[30][39],
reservoir_weight[30][40],
reservoir_weight[30][41],
reservoir_weight[30][42],
reservoir_weight[30][43],
reservoir_weight[30][44],
reservoir_weight[30][45],
reservoir_weight[30][46],
reservoir_weight[30][47],
reservoir_weight[30][48],
reservoir_weight[30][49],
reservoir_weight[30][50],
reservoir_weight[30][51],
reservoir_weight[30][52],
reservoir_weight[30][53],
reservoir_weight[30][54],
reservoir_weight[30][55],
reservoir_weight[30][56],
reservoir_weight[30][57],
reservoir_weight[30][58],
reservoir_weight[30][59],
reservoir_weight[30][60],
reservoir_weight[30][61],
reservoir_weight[30][62],
reservoir_weight[30][63],
reservoir_weight[30][64],
reservoir_weight[30][65],
reservoir_weight[30][66],
reservoir_weight[30][67],
reservoir_weight[30][68],
reservoir_weight[30][69],
reservoir_weight[30][70],
reservoir_weight[30][71],
reservoir_weight[30][72],
reservoir_weight[30][73],
reservoir_weight[30][74],
reservoir_weight[30][75],
reservoir_weight[30][76],
reservoir_weight[30][77],
reservoir_weight[30][78],
reservoir_weight[30][79],
reservoir_weight[30][80],
reservoir_weight[30][81],
reservoir_weight[30][82],
reservoir_weight[30][83],
reservoir_weight[30][84],
reservoir_weight[30][85],
reservoir_weight[30][86],
reservoir_weight[30][87],
reservoir_weight[30][88],
reservoir_weight[30][89],
reservoir_weight[30][90],
reservoir_weight[30][91],
reservoir_weight[30][92],
reservoir_weight[30][93],
reservoir_weight[30][94],
reservoir_weight[30][95],
reservoir_weight[30][96],
reservoir_weight[30][97],
reservoir_weight[30][98],
reservoir_weight[30][99],
reservoir_weight[30][100],
reservoir_weight[30][101],
reservoir_weight[30][102],
reservoir_weight[30][103],
reservoir_weight[30][104],
reservoir_weight[30][105],
reservoir_weight[30][106],
reservoir_weight[30][107],
reservoir_weight[30][108],
reservoir_weight[30][109],
reservoir_weight[30][110],
reservoir_weight[30][111],
reservoir_weight[30][112],
reservoir_weight[30][113],
reservoir_weight[30][114],
reservoir_weight[30][115],
reservoir_weight[30][116],
reservoir_weight[30][117],
reservoir_weight[30][118],
reservoir_weight[30][119],
reservoir_weight[30][120],
reservoir_weight[30][121],
reservoir_weight[30][122],
reservoir_weight[30][123],
reservoir_weight[30][124],
reservoir_weight[30][125],
reservoir_weight[30][126],
reservoir_weight[30][127],
reservoir_weight[30][128],
reservoir_weight[30][129],
reservoir_weight[30][130],
reservoir_weight[30][131],
reservoir_weight[30][132],
reservoir_weight[30][133],
reservoir_weight[30][134],
reservoir_weight[30][135],
reservoir_weight[30][136],
reservoir_weight[30][137],
reservoir_weight[30][138],
reservoir_weight[30][139],
reservoir_weight[30][140],
reservoir_weight[30][141],
reservoir_weight[30][142],
reservoir_weight[30][143],
reservoir_weight[30][144],
reservoir_weight[30][145],
reservoir_weight[30][146],
reservoir_weight[30][147],
reservoir_weight[30][148],
reservoir_weight[30][149],
reservoir_weight[30][150],
reservoir_weight[30][151],
reservoir_weight[30][152],
reservoir_weight[30][153],
reservoir_weight[30][154],
reservoir_weight[30][155],
reservoir_weight[30][156],
reservoir_weight[30][157],
reservoir_weight[30][158],
reservoir_weight[30][159],
reservoir_weight[30][160],
reservoir_weight[30][161],
reservoir_weight[30][162],
reservoir_weight[30][163],
reservoir_weight[30][164],
reservoir_weight[30][165],
reservoir_weight[30][166],
reservoir_weight[30][167],
reservoir_weight[30][168],
reservoir_weight[30][169],
reservoir_weight[30][170],
reservoir_weight[30][171],
reservoir_weight[30][172],
reservoir_weight[30][173],
reservoir_weight[30][174],
reservoir_weight[30][175],
reservoir_weight[30][176],
reservoir_weight[30][177],
reservoir_weight[30][178],
reservoir_weight[30][179],
reservoir_weight[30][180],
reservoir_weight[30][181],
reservoir_weight[30][182],
reservoir_weight[30][183],
reservoir_weight[30][184],
reservoir_weight[30][185],
reservoir_weight[30][186],
reservoir_weight[30][187],
reservoir_weight[30][188],
reservoir_weight[30][189],
reservoir_weight[30][190],
reservoir_weight[30][191],
reservoir_weight[30][192],
reservoir_weight[30][193],
reservoir_weight[30][194],
reservoir_weight[30][195],
reservoir_weight[30][196],
reservoir_weight[30][197],
reservoir_weight[30][198],
reservoir_weight[30][199]
},
{reservoir_weight[31][0],
reservoir_weight[31][1],
reservoir_weight[31][2],
reservoir_weight[31][3],
reservoir_weight[31][4],
reservoir_weight[31][5],
reservoir_weight[31][6],
reservoir_weight[31][7],
reservoir_weight[31][8],
reservoir_weight[31][9],
reservoir_weight[31][10],
reservoir_weight[31][11],
reservoir_weight[31][12],
reservoir_weight[31][13],
reservoir_weight[31][14],
reservoir_weight[31][15],
reservoir_weight[31][16],
reservoir_weight[31][17],
reservoir_weight[31][18],
reservoir_weight[31][19],
reservoir_weight[31][20],
reservoir_weight[31][21],
reservoir_weight[31][22],
reservoir_weight[31][23],
reservoir_weight[31][24],
reservoir_weight[31][25],
reservoir_weight[31][26],
reservoir_weight[31][27],
reservoir_weight[31][28],
reservoir_weight[31][29],
reservoir_weight[31][30],
reservoir_weight[31][31],
reservoir_weight[31][32],
reservoir_weight[31][33],
reservoir_weight[31][34],
reservoir_weight[31][35],
reservoir_weight[31][36],
reservoir_weight[31][37],
reservoir_weight[31][38],
reservoir_weight[31][39],
reservoir_weight[31][40],
reservoir_weight[31][41],
reservoir_weight[31][42],
reservoir_weight[31][43],
reservoir_weight[31][44],
reservoir_weight[31][45],
reservoir_weight[31][46],
reservoir_weight[31][47],
reservoir_weight[31][48],
reservoir_weight[31][49],
reservoir_weight[31][50],
reservoir_weight[31][51],
reservoir_weight[31][52],
reservoir_weight[31][53],
reservoir_weight[31][54],
reservoir_weight[31][55],
reservoir_weight[31][56],
reservoir_weight[31][57],
reservoir_weight[31][58],
reservoir_weight[31][59],
reservoir_weight[31][60],
reservoir_weight[31][61],
reservoir_weight[31][62],
reservoir_weight[31][63],
reservoir_weight[31][64],
reservoir_weight[31][65],
reservoir_weight[31][66],
reservoir_weight[31][67],
reservoir_weight[31][68],
reservoir_weight[31][69],
reservoir_weight[31][70],
reservoir_weight[31][71],
reservoir_weight[31][72],
reservoir_weight[31][73],
reservoir_weight[31][74],
reservoir_weight[31][75],
reservoir_weight[31][76],
reservoir_weight[31][77],
reservoir_weight[31][78],
reservoir_weight[31][79],
reservoir_weight[31][80],
reservoir_weight[31][81],
reservoir_weight[31][82],
reservoir_weight[31][83],
reservoir_weight[31][84],
reservoir_weight[31][85],
reservoir_weight[31][86],
reservoir_weight[31][87],
reservoir_weight[31][88],
reservoir_weight[31][89],
reservoir_weight[31][90],
reservoir_weight[31][91],
reservoir_weight[31][92],
reservoir_weight[31][93],
reservoir_weight[31][94],
reservoir_weight[31][95],
reservoir_weight[31][96],
reservoir_weight[31][97],
reservoir_weight[31][98],
reservoir_weight[31][99],
reservoir_weight[31][100],
reservoir_weight[31][101],
reservoir_weight[31][102],
reservoir_weight[31][103],
reservoir_weight[31][104],
reservoir_weight[31][105],
reservoir_weight[31][106],
reservoir_weight[31][107],
reservoir_weight[31][108],
reservoir_weight[31][109],
reservoir_weight[31][110],
reservoir_weight[31][111],
reservoir_weight[31][112],
reservoir_weight[31][113],
reservoir_weight[31][114],
reservoir_weight[31][115],
reservoir_weight[31][116],
reservoir_weight[31][117],
reservoir_weight[31][118],
reservoir_weight[31][119],
reservoir_weight[31][120],
reservoir_weight[31][121],
reservoir_weight[31][122],
reservoir_weight[31][123],
reservoir_weight[31][124],
reservoir_weight[31][125],
reservoir_weight[31][126],
reservoir_weight[31][127],
reservoir_weight[31][128],
reservoir_weight[31][129],
reservoir_weight[31][130],
reservoir_weight[31][131],
reservoir_weight[31][132],
reservoir_weight[31][133],
reservoir_weight[31][134],
reservoir_weight[31][135],
reservoir_weight[31][136],
reservoir_weight[31][137],
reservoir_weight[31][138],
reservoir_weight[31][139],
reservoir_weight[31][140],
reservoir_weight[31][141],
reservoir_weight[31][142],
reservoir_weight[31][143],
reservoir_weight[31][144],
reservoir_weight[31][145],
reservoir_weight[31][146],
reservoir_weight[31][147],
reservoir_weight[31][148],
reservoir_weight[31][149],
reservoir_weight[31][150],
reservoir_weight[31][151],
reservoir_weight[31][152],
reservoir_weight[31][153],
reservoir_weight[31][154],
reservoir_weight[31][155],
reservoir_weight[31][156],
reservoir_weight[31][157],
reservoir_weight[31][158],
reservoir_weight[31][159],
reservoir_weight[31][160],
reservoir_weight[31][161],
reservoir_weight[31][162],
reservoir_weight[31][163],
reservoir_weight[31][164],
reservoir_weight[31][165],
reservoir_weight[31][166],
reservoir_weight[31][167],
reservoir_weight[31][168],
reservoir_weight[31][169],
reservoir_weight[31][170],
reservoir_weight[31][171],
reservoir_weight[31][172],
reservoir_weight[31][173],
reservoir_weight[31][174],
reservoir_weight[31][175],
reservoir_weight[31][176],
reservoir_weight[31][177],
reservoir_weight[31][178],
reservoir_weight[31][179],
reservoir_weight[31][180],
reservoir_weight[31][181],
reservoir_weight[31][182],
reservoir_weight[31][183],
reservoir_weight[31][184],
reservoir_weight[31][185],
reservoir_weight[31][186],
reservoir_weight[31][187],
reservoir_weight[31][188],
reservoir_weight[31][189],
reservoir_weight[31][190],
reservoir_weight[31][191],
reservoir_weight[31][192],
reservoir_weight[31][193],
reservoir_weight[31][194],
reservoir_weight[31][195],
reservoir_weight[31][196],
reservoir_weight[31][197],
reservoir_weight[31][198],
reservoir_weight[31][199]
},
{reservoir_weight[32][0],
reservoir_weight[32][1],
reservoir_weight[32][2],
reservoir_weight[32][3],
reservoir_weight[32][4],
reservoir_weight[32][5],
reservoir_weight[32][6],
reservoir_weight[32][7],
reservoir_weight[32][8],
reservoir_weight[32][9],
reservoir_weight[32][10],
reservoir_weight[32][11],
reservoir_weight[32][12],
reservoir_weight[32][13],
reservoir_weight[32][14],
reservoir_weight[32][15],
reservoir_weight[32][16],
reservoir_weight[32][17],
reservoir_weight[32][18],
reservoir_weight[32][19],
reservoir_weight[32][20],
reservoir_weight[32][21],
reservoir_weight[32][22],
reservoir_weight[32][23],
reservoir_weight[32][24],
reservoir_weight[32][25],
reservoir_weight[32][26],
reservoir_weight[32][27],
reservoir_weight[32][28],
reservoir_weight[32][29],
reservoir_weight[32][30],
reservoir_weight[32][31],
reservoir_weight[32][32],
reservoir_weight[32][33],
reservoir_weight[32][34],
reservoir_weight[32][35],
reservoir_weight[32][36],
reservoir_weight[32][37],
reservoir_weight[32][38],
reservoir_weight[32][39],
reservoir_weight[32][40],
reservoir_weight[32][41],
reservoir_weight[32][42],
reservoir_weight[32][43],
reservoir_weight[32][44],
reservoir_weight[32][45],
reservoir_weight[32][46],
reservoir_weight[32][47],
reservoir_weight[32][48],
reservoir_weight[32][49],
reservoir_weight[32][50],
reservoir_weight[32][51],
reservoir_weight[32][52],
reservoir_weight[32][53],
reservoir_weight[32][54],
reservoir_weight[32][55],
reservoir_weight[32][56],
reservoir_weight[32][57],
reservoir_weight[32][58],
reservoir_weight[32][59],
reservoir_weight[32][60],
reservoir_weight[32][61],
reservoir_weight[32][62],
reservoir_weight[32][63],
reservoir_weight[32][64],
reservoir_weight[32][65],
reservoir_weight[32][66],
reservoir_weight[32][67],
reservoir_weight[32][68],
reservoir_weight[32][69],
reservoir_weight[32][70],
reservoir_weight[32][71],
reservoir_weight[32][72],
reservoir_weight[32][73],
reservoir_weight[32][74],
reservoir_weight[32][75],
reservoir_weight[32][76],
reservoir_weight[32][77],
reservoir_weight[32][78],
reservoir_weight[32][79],
reservoir_weight[32][80],
reservoir_weight[32][81],
reservoir_weight[32][82],
reservoir_weight[32][83],
reservoir_weight[32][84],
reservoir_weight[32][85],
reservoir_weight[32][86],
reservoir_weight[32][87],
reservoir_weight[32][88],
reservoir_weight[32][89],
reservoir_weight[32][90],
reservoir_weight[32][91],
reservoir_weight[32][92],
reservoir_weight[32][93],
reservoir_weight[32][94],
reservoir_weight[32][95],
reservoir_weight[32][96],
reservoir_weight[32][97],
reservoir_weight[32][98],
reservoir_weight[32][99],
reservoir_weight[32][100],
reservoir_weight[32][101],
reservoir_weight[32][102],
reservoir_weight[32][103],
reservoir_weight[32][104],
reservoir_weight[32][105],
reservoir_weight[32][106],
reservoir_weight[32][107],
reservoir_weight[32][108],
reservoir_weight[32][109],
reservoir_weight[32][110],
reservoir_weight[32][111],
reservoir_weight[32][112],
reservoir_weight[32][113],
reservoir_weight[32][114],
reservoir_weight[32][115],
reservoir_weight[32][116],
reservoir_weight[32][117],
reservoir_weight[32][118],
reservoir_weight[32][119],
reservoir_weight[32][120],
reservoir_weight[32][121],
reservoir_weight[32][122],
reservoir_weight[32][123],
reservoir_weight[32][124],
reservoir_weight[32][125],
reservoir_weight[32][126],
reservoir_weight[32][127],
reservoir_weight[32][128],
reservoir_weight[32][129],
reservoir_weight[32][130],
reservoir_weight[32][131],
reservoir_weight[32][132],
reservoir_weight[32][133],
reservoir_weight[32][134],
reservoir_weight[32][135],
reservoir_weight[32][136],
reservoir_weight[32][137],
reservoir_weight[32][138],
reservoir_weight[32][139],
reservoir_weight[32][140],
reservoir_weight[32][141],
reservoir_weight[32][142],
reservoir_weight[32][143],
reservoir_weight[32][144],
reservoir_weight[32][145],
reservoir_weight[32][146],
reservoir_weight[32][147],
reservoir_weight[32][148],
reservoir_weight[32][149],
reservoir_weight[32][150],
reservoir_weight[32][151],
reservoir_weight[32][152],
reservoir_weight[32][153],
reservoir_weight[32][154],
reservoir_weight[32][155],
reservoir_weight[32][156],
reservoir_weight[32][157],
reservoir_weight[32][158],
reservoir_weight[32][159],
reservoir_weight[32][160],
reservoir_weight[32][161],
reservoir_weight[32][162],
reservoir_weight[32][163],
reservoir_weight[32][164],
reservoir_weight[32][165],
reservoir_weight[32][166],
reservoir_weight[32][167],
reservoir_weight[32][168],
reservoir_weight[32][169],
reservoir_weight[32][170],
reservoir_weight[32][171],
reservoir_weight[32][172],
reservoir_weight[32][173],
reservoir_weight[32][174],
reservoir_weight[32][175],
reservoir_weight[32][176],
reservoir_weight[32][177],
reservoir_weight[32][178],
reservoir_weight[32][179],
reservoir_weight[32][180],
reservoir_weight[32][181],
reservoir_weight[32][182],
reservoir_weight[32][183],
reservoir_weight[32][184],
reservoir_weight[32][185],
reservoir_weight[32][186],
reservoir_weight[32][187],
reservoir_weight[32][188],
reservoir_weight[32][189],
reservoir_weight[32][190],
reservoir_weight[32][191],
reservoir_weight[32][192],
reservoir_weight[32][193],
reservoir_weight[32][194],
reservoir_weight[32][195],
reservoir_weight[32][196],
reservoir_weight[32][197],
reservoir_weight[32][198],
reservoir_weight[32][199]
},
{reservoir_weight[33][0],
reservoir_weight[33][1],
reservoir_weight[33][2],
reservoir_weight[33][3],
reservoir_weight[33][4],
reservoir_weight[33][5],
reservoir_weight[33][6],
reservoir_weight[33][7],
reservoir_weight[33][8],
reservoir_weight[33][9],
reservoir_weight[33][10],
reservoir_weight[33][11],
reservoir_weight[33][12],
reservoir_weight[33][13],
reservoir_weight[33][14],
reservoir_weight[33][15],
reservoir_weight[33][16],
reservoir_weight[33][17],
reservoir_weight[33][18],
reservoir_weight[33][19],
reservoir_weight[33][20],
reservoir_weight[33][21],
reservoir_weight[33][22],
reservoir_weight[33][23],
reservoir_weight[33][24],
reservoir_weight[33][25],
reservoir_weight[33][26],
reservoir_weight[33][27],
reservoir_weight[33][28],
reservoir_weight[33][29],
reservoir_weight[33][30],
reservoir_weight[33][31],
reservoir_weight[33][32],
reservoir_weight[33][33],
reservoir_weight[33][34],
reservoir_weight[33][35],
reservoir_weight[33][36],
reservoir_weight[33][37],
reservoir_weight[33][38],
reservoir_weight[33][39],
reservoir_weight[33][40],
reservoir_weight[33][41],
reservoir_weight[33][42],
reservoir_weight[33][43],
reservoir_weight[33][44],
reservoir_weight[33][45],
reservoir_weight[33][46],
reservoir_weight[33][47],
reservoir_weight[33][48],
reservoir_weight[33][49],
reservoir_weight[33][50],
reservoir_weight[33][51],
reservoir_weight[33][52],
reservoir_weight[33][53],
reservoir_weight[33][54],
reservoir_weight[33][55],
reservoir_weight[33][56],
reservoir_weight[33][57],
reservoir_weight[33][58],
reservoir_weight[33][59],
reservoir_weight[33][60],
reservoir_weight[33][61],
reservoir_weight[33][62],
reservoir_weight[33][63],
reservoir_weight[33][64],
reservoir_weight[33][65],
reservoir_weight[33][66],
reservoir_weight[33][67],
reservoir_weight[33][68],
reservoir_weight[33][69],
reservoir_weight[33][70],
reservoir_weight[33][71],
reservoir_weight[33][72],
reservoir_weight[33][73],
reservoir_weight[33][74],
reservoir_weight[33][75],
reservoir_weight[33][76],
reservoir_weight[33][77],
reservoir_weight[33][78],
reservoir_weight[33][79],
reservoir_weight[33][80],
reservoir_weight[33][81],
reservoir_weight[33][82],
reservoir_weight[33][83],
reservoir_weight[33][84],
reservoir_weight[33][85],
reservoir_weight[33][86],
reservoir_weight[33][87],
reservoir_weight[33][88],
reservoir_weight[33][89],
reservoir_weight[33][90],
reservoir_weight[33][91],
reservoir_weight[33][92],
reservoir_weight[33][93],
reservoir_weight[33][94],
reservoir_weight[33][95],
reservoir_weight[33][96],
reservoir_weight[33][97],
reservoir_weight[33][98],
reservoir_weight[33][99],
reservoir_weight[33][100],
reservoir_weight[33][101],
reservoir_weight[33][102],
reservoir_weight[33][103],
reservoir_weight[33][104],
reservoir_weight[33][105],
reservoir_weight[33][106],
reservoir_weight[33][107],
reservoir_weight[33][108],
reservoir_weight[33][109],
reservoir_weight[33][110],
reservoir_weight[33][111],
reservoir_weight[33][112],
reservoir_weight[33][113],
reservoir_weight[33][114],
reservoir_weight[33][115],
reservoir_weight[33][116],
reservoir_weight[33][117],
reservoir_weight[33][118],
reservoir_weight[33][119],
reservoir_weight[33][120],
reservoir_weight[33][121],
reservoir_weight[33][122],
reservoir_weight[33][123],
reservoir_weight[33][124],
reservoir_weight[33][125],
reservoir_weight[33][126],
reservoir_weight[33][127],
reservoir_weight[33][128],
reservoir_weight[33][129],
reservoir_weight[33][130],
reservoir_weight[33][131],
reservoir_weight[33][132],
reservoir_weight[33][133],
reservoir_weight[33][134],
reservoir_weight[33][135],
reservoir_weight[33][136],
reservoir_weight[33][137],
reservoir_weight[33][138],
reservoir_weight[33][139],
reservoir_weight[33][140],
reservoir_weight[33][141],
reservoir_weight[33][142],
reservoir_weight[33][143],
reservoir_weight[33][144],
reservoir_weight[33][145],
reservoir_weight[33][146],
reservoir_weight[33][147],
reservoir_weight[33][148],
reservoir_weight[33][149],
reservoir_weight[33][150],
reservoir_weight[33][151],
reservoir_weight[33][152],
reservoir_weight[33][153],
reservoir_weight[33][154],
reservoir_weight[33][155],
reservoir_weight[33][156],
reservoir_weight[33][157],
reservoir_weight[33][158],
reservoir_weight[33][159],
reservoir_weight[33][160],
reservoir_weight[33][161],
reservoir_weight[33][162],
reservoir_weight[33][163],
reservoir_weight[33][164],
reservoir_weight[33][165],
reservoir_weight[33][166],
reservoir_weight[33][167],
reservoir_weight[33][168],
reservoir_weight[33][169],
reservoir_weight[33][170],
reservoir_weight[33][171],
reservoir_weight[33][172],
reservoir_weight[33][173],
reservoir_weight[33][174],
reservoir_weight[33][175],
reservoir_weight[33][176],
reservoir_weight[33][177],
reservoir_weight[33][178],
reservoir_weight[33][179],
reservoir_weight[33][180],
reservoir_weight[33][181],
reservoir_weight[33][182],
reservoir_weight[33][183],
reservoir_weight[33][184],
reservoir_weight[33][185],
reservoir_weight[33][186],
reservoir_weight[33][187],
reservoir_weight[33][188],
reservoir_weight[33][189],
reservoir_weight[33][190],
reservoir_weight[33][191],
reservoir_weight[33][192],
reservoir_weight[33][193],
reservoir_weight[33][194],
reservoir_weight[33][195],
reservoir_weight[33][196],
reservoir_weight[33][197],
reservoir_weight[33][198],
reservoir_weight[33][199]
},
{reservoir_weight[34][0],
reservoir_weight[34][1],
reservoir_weight[34][2],
reservoir_weight[34][3],
reservoir_weight[34][4],
reservoir_weight[34][5],
reservoir_weight[34][6],
reservoir_weight[34][7],
reservoir_weight[34][8],
reservoir_weight[34][9],
reservoir_weight[34][10],
reservoir_weight[34][11],
reservoir_weight[34][12],
reservoir_weight[34][13],
reservoir_weight[34][14],
reservoir_weight[34][15],
reservoir_weight[34][16],
reservoir_weight[34][17],
reservoir_weight[34][18],
reservoir_weight[34][19],
reservoir_weight[34][20],
reservoir_weight[34][21],
reservoir_weight[34][22],
reservoir_weight[34][23],
reservoir_weight[34][24],
reservoir_weight[34][25],
reservoir_weight[34][26],
reservoir_weight[34][27],
reservoir_weight[34][28],
reservoir_weight[34][29],
reservoir_weight[34][30],
reservoir_weight[34][31],
reservoir_weight[34][32],
reservoir_weight[34][33],
reservoir_weight[34][34],
reservoir_weight[34][35],
reservoir_weight[34][36],
reservoir_weight[34][37],
reservoir_weight[34][38],
reservoir_weight[34][39],
reservoir_weight[34][40],
reservoir_weight[34][41],
reservoir_weight[34][42],
reservoir_weight[34][43],
reservoir_weight[34][44],
reservoir_weight[34][45],
reservoir_weight[34][46],
reservoir_weight[34][47],
reservoir_weight[34][48],
reservoir_weight[34][49],
reservoir_weight[34][50],
reservoir_weight[34][51],
reservoir_weight[34][52],
reservoir_weight[34][53],
reservoir_weight[34][54],
reservoir_weight[34][55],
reservoir_weight[34][56],
reservoir_weight[34][57],
reservoir_weight[34][58],
reservoir_weight[34][59],
reservoir_weight[34][60],
reservoir_weight[34][61],
reservoir_weight[34][62],
reservoir_weight[34][63],
reservoir_weight[34][64],
reservoir_weight[34][65],
reservoir_weight[34][66],
reservoir_weight[34][67],
reservoir_weight[34][68],
reservoir_weight[34][69],
reservoir_weight[34][70],
reservoir_weight[34][71],
reservoir_weight[34][72],
reservoir_weight[34][73],
reservoir_weight[34][74],
reservoir_weight[34][75],
reservoir_weight[34][76],
reservoir_weight[34][77],
reservoir_weight[34][78],
reservoir_weight[34][79],
reservoir_weight[34][80],
reservoir_weight[34][81],
reservoir_weight[34][82],
reservoir_weight[34][83],
reservoir_weight[34][84],
reservoir_weight[34][85],
reservoir_weight[34][86],
reservoir_weight[34][87],
reservoir_weight[34][88],
reservoir_weight[34][89],
reservoir_weight[34][90],
reservoir_weight[34][91],
reservoir_weight[34][92],
reservoir_weight[34][93],
reservoir_weight[34][94],
reservoir_weight[34][95],
reservoir_weight[34][96],
reservoir_weight[34][97],
reservoir_weight[34][98],
reservoir_weight[34][99],
reservoir_weight[34][100],
reservoir_weight[34][101],
reservoir_weight[34][102],
reservoir_weight[34][103],
reservoir_weight[34][104],
reservoir_weight[34][105],
reservoir_weight[34][106],
reservoir_weight[34][107],
reservoir_weight[34][108],
reservoir_weight[34][109],
reservoir_weight[34][110],
reservoir_weight[34][111],
reservoir_weight[34][112],
reservoir_weight[34][113],
reservoir_weight[34][114],
reservoir_weight[34][115],
reservoir_weight[34][116],
reservoir_weight[34][117],
reservoir_weight[34][118],
reservoir_weight[34][119],
reservoir_weight[34][120],
reservoir_weight[34][121],
reservoir_weight[34][122],
reservoir_weight[34][123],
reservoir_weight[34][124],
reservoir_weight[34][125],
reservoir_weight[34][126],
reservoir_weight[34][127],
reservoir_weight[34][128],
reservoir_weight[34][129],
reservoir_weight[34][130],
reservoir_weight[34][131],
reservoir_weight[34][132],
reservoir_weight[34][133],
reservoir_weight[34][134],
reservoir_weight[34][135],
reservoir_weight[34][136],
reservoir_weight[34][137],
reservoir_weight[34][138],
reservoir_weight[34][139],
reservoir_weight[34][140],
reservoir_weight[34][141],
reservoir_weight[34][142],
reservoir_weight[34][143],
reservoir_weight[34][144],
reservoir_weight[34][145],
reservoir_weight[34][146],
reservoir_weight[34][147],
reservoir_weight[34][148],
reservoir_weight[34][149],
reservoir_weight[34][150],
reservoir_weight[34][151],
reservoir_weight[34][152],
reservoir_weight[34][153],
reservoir_weight[34][154],
reservoir_weight[34][155],
reservoir_weight[34][156],
reservoir_weight[34][157],
reservoir_weight[34][158],
reservoir_weight[34][159],
reservoir_weight[34][160],
reservoir_weight[34][161],
reservoir_weight[34][162],
reservoir_weight[34][163],
reservoir_weight[34][164],
reservoir_weight[34][165],
reservoir_weight[34][166],
reservoir_weight[34][167],
reservoir_weight[34][168],
reservoir_weight[34][169],
reservoir_weight[34][170],
reservoir_weight[34][171],
reservoir_weight[34][172],
reservoir_weight[34][173],
reservoir_weight[34][174],
reservoir_weight[34][175],
reservoir_weight[34][176],
reservoir_weight[34][177],
reservoir_weight[34][178],
reservoir_weight[34][179],
reservoir_weight[34][180],
reservoir_weight[34][181],
reservoir_weight[34][182],
reservoir_weight[34][183],
reservoir_weight[34][184],
reservoir_weight[34][185],
reservoir_weight[34][186],
reservoir_weight[34][187],
reservoir_weight[34][188],
reservoir_weight[34][189],
reservoir_weight[34][190],
reservoir_weight[34][191],
reservoir_weight[34][192],
reservoir_weight[34][193],
reservoir_weight[34][194],
reservoir_weight[34][195],
reservoir_weight[34][196],
reservoir_weight[34][197],
reservoir_weight[34][198],
reservoir_weight[34][199]
},
{reservoir_weight[35][0],
reservoir_weight[35][1],
reservoir_weight[35][2],
reservoir_weight[35][3],
reservoir_weight[35][4],
reservoir_weight[35][5],
reservoir_weight[35][6],
reservoir_weight[35][7],
reservoir_weight[35][8],
reservoir_weight[35][9],
reservoir_weight[35][10],
reservoir_weight[35][11],
reservoir_weight[35][12],
reservoir_weight[35][13],
reservoir_weight[35][14],
reservoir_weight[35][15],
reservoir_weight[35][16],
reservoir_weight[35][17],
reservoir_weight[35][18],
reservoir_weight[35][19],
reservoir_weight[35][20],
reservoir_weight[35][21],
reservoir_weight[35][22],
reservoir_weight[35][23],
reservoir_weight[35][24],
reservoir_weight[35][25],
reservoir_weight[35][26],
reservoir_weight[35][27],
reservoir_weight[35][28],
reservoir_weight[35][29],
reservoir_weight[35][30],
reservoir_weight[35][31],
reservoir_weight[35][32],
reservoir_weight[35][33],
reservoir_weight[35][34],
reservoir_weight[35][35],
reservoir_weight[35][36],
reservoir_weight[35][37],
reservoir_weight[35][38],
reservoir_weight[35][39],
reservoir_weight[35][40],
reservoir_weight[35][41],
reservoir_weight[35][42],
reservoir_weight[35][43],
reservoir_weight[35][44],
reservoir_weight[35][45],
reservoir_weight[35][46],
reservoir_weight[35][47],
reservoir_weight[35][48],
reservoir_weight[35][49],
reservoir_weight[35][50],
reservoir_weight[35][51],
reservoir_weight[35][52],
reservoir_weight[35][53],
reservoir_weight[35][54],
reservoir_weight[35][55],
reservoir_weight[35][56],
reservoir_weight[35][57],
reservoir_weight[35][58],
reservoir_weight[35][59],
reservoir_weight[35][60],
reservoir_weight[35][61],
reservoir_weight[35][62],
reservoir_weight[35][63],
reservoir_weight[35][64],
reservoir_weight[35][65],
reservoir_weight[35][66],
reservoir_weight[35][67],
reservoir_weight[35][68],
reservoir_weight[35][69],
reservoir_weight[35][70],
reservoir_weight[35][71],
reservoir_weight[35][72],
reservoir_weight[35][73],
reservoir_weight[35][74],
reservoir_weight[35][75],
reservoir_weight[35][76],
reservoir_weight[35][77],
reservoir_weight[35][78],
reservoir_weight[35][79],
reservoir_weight[35][80],
reservoir_weight[35][81],
reservoir_weight[35][82],
reservoir_weight[35][83],
reservoir_weight[35][84],
reservoir_weight[35][85],
reservoir_weight[35][86],
reservoir_weight[35][87],
reservoir_weight[35][88],
reservoir_weight[35][89],
reservoir_weight[35][90],
reservoir_weight[35][91],
reservoir_weight[35][92],
reservoir_weight[35][93],
reservoir_weight[35][94],
reservoir_weight[35][95],
reservoir_weight[35][96],
reservoir_weight[35][97],
reservoir_weight[35][98],
reservoir_weight[35][99],
reservoir_weight[35][100],
reservoir_weight[35][101],
reservoir_weight[35][102],
reservoir_weight[35][103],
reservoir_weight[35][104],
reservoir_weight[35][105],
reservoir_weight[35][106],
reservoir_weight[35][107],
reservoir_weight[35][108],
reservoir_weight[35][109],
reservoir_weight[35][110],
reservoir_weight[35][111],
reservoir_weight[35][112],
reservoir_weight[35][113],
reservoir_weight[35][114],
reservoir_weight[35][115],
reservoir_weight[35][116],
reservoir_weight[35][117],
reservoir_weight[35][118],
reservoir_weight[35][119],
reservoir_weight[35][120],
reservoir_weight[35][121],
reservoir_weight[35][122],
reservoir_weight[35][123],
reservoir_weight[35][124],
reservoir_weight[35][125],
reservoir_weight[35][126],
reservoir_weight[35][127],
reservoir_weight[35][128],
reservoir_weight[35][129],
reservoir_weight[35][130],
reservoir_weight[35][131],
reservoir_weight[35][132],
reservoir_weight[35][133],
reservoir_weight[35][134],
reservoir_weight[35][135],
reservoir_weight[35][136],
reservoir_weight[35][137],
reservoir_weight[35][138],
reservoir_weight[35][139],
reservoir_weight[35][140],
reservoir_weight[35][141],
reservoir_weight[35][142],
reservoir_weight[35][143],
reservoir_weight[35][144],
reservoir_weight[35][145],
reservoir_weight[35][146],
reservoir_weight[35][147],
reservoir_weight[35][148],
reservoir_weight[35][149],
reservoir_weight[35][150],
reservoir_weight[35][151],
reservoir_weight[35][152],
reservoir_weight[35][153],
reservoir_weight[35][154],
reservoir_weight[35][155],
reservoir_weight[35][156],
reservoir_weight[35][157],
reservoir_weight[35][158],
reservoir_weight[35][159],
reservoir_weight[35][160],
reservoir_weight[35][161],
reservoir_weight[35][162],
reservoir_weight[35][163],
reservoir_weight[35][164],
reservoir_weight[35][165],
reservoir_weight[35][166],
reservoir_weight[35][167],
reservoir_weight[35][168],
reservoir_weight[35][169],
reservoir_weight[35][170],
reservoir_weight[35][171],
reservoir_weight[35][172],
reservoir_weight[35][173],
reservoir_weight[35][174],
reservoir_weight[35][175],
reservoir_weight[35][176],
reservoir_weight[35][177],
reservoir_weight[35][178],
reservoir_weight[35][179],
reservoir_weight[35][180],
reservoir_weight[35][181],
reservoir_weight[35][182],
reservoir_weight[35][183],
reservoir_weight[35][184],
reservoir_weight[35][185],
reservoir_weight[35][186],
reservoir_weight[35][187],
reservoir_weight[35][188],
reservoir_weight[35][189],
reservoir_weight[35][190],
reservoir_weight[35][191],
reservoir_weight[35][192],
reservoir_weight[35][193],
reservoir_weight[35][194],
reservoir_weight[35][195],
reservoir_weight[35][196],
reservoir_weight[35][197],
reservoir_weight[35][198],
reservoir_weight[35][199]
},
{reservoir_weight[36][0],
reservoir_weight[36][1],
reservoir_weight[36][2],
reservoir_weight[36][3],
reservoir_weight[36][4],
reservoir_weight[36][5],
reservoir_weight[36][6],
reservoir_weight[36][7],
reservoir_weight[36][8],
reservoir_weight[36][9],
reservoir_weight[36][10],
reservoir_weight[36][11],
reservoir_weight[36][12],
reservoir_weight[36][13],
reservoir_weight[36][14],
reservoir_weight[36][15],
reservoir_weight[36][16],
reservoir_weight[36][17],
reservoir_weight[36][18],
reservoir_weight[36][19],
reservoir_weight[36][20],
reservoir_weight[36][21],
reservoir_weight[36][22],
reservoir_weight[36][23],
reservoir_weight[36][24],
reservoir_weight[36][25],
reservoir_weight[36][26],
reservoir_weight[36][27],
reservoir_weight[36][28],
reservoir_weight[36][29],
reservoir_weight[36][30],
reservoir_weight[36][31],
reservoir_weight[36][32],
reservoir_weight[36][33],
reservoir_weight[36][34],
reservoir_weight[36][35],
reservoir_weight[36][36],
reservoir_weight[36][37],
reservoir_weight[36][38],
reservoir_weight[36][39],
reservoir_weight[36][40],
reservoir_weight[36][41],
reservoir_weight[36][42],
reservoir_weight[36][43],
reservoir_weight[36][44],
reservoir_weight[36][45],
reservoir_weight[36][46],
reservoir_weight[36][47],
reservoir_weight[36][48],
reservoir_weight[36][49],
reservoir_weight[36][50],
reservoir_weight[36][51],
reservoir_weight[36][52],
reservoir_weight[36][53],
reservoir_weight[36][54],
reservoir_weight[36][55],
reservoir_weight[36][56],
reservoir_weight[36][57],
reservoir_weight[36][58],
reservoir_weight[36][59],
reservoir_weight[36][60],
reservoir_weight[36][61],
reservoir_weight[36][62],
reservoir_weight[36][63],
reservoir_weight[36][64],
reservoir_weight[36][65],
reservoir_weight[36][66],
reservoir_weight[36][67],
reservoir_weight[36][68],
reservoir_weight[36][69],
reservoir_weight[36][70],
reservoir_weight[36][71],
reservoir_weight[36][72],
reservoir_weight[36][73],
reservoir_weight[36][74],
reservoir_weight[36][75],
reservoir_weight[36][76],
reservoir_weight[36][77],
reservoir_weight[36][78],
reservoir_weight[36][79],
reservoir_weight[36][80],
reservoir_weight[36][81],
reservoir_weight[36][82],
reservoir_weight[36][83],
reservoir_weight[36][84],
reservoir_weight[36][85],
reservoir_weight[36][86],
reservoir_weight[36][87],
reservoir_weight[36][88],
reservoir_weight[36][89],
reservoir_weight[36][90],
reservoir_weight[36][91],
reservoir_weight[36][92],
reservoir_weight[36][93],
reservoir_weight[36][94],
reservoir_weight[36][95],
reservoir_weight[36][96],
reservoir_weight[36][97],
reservoir_weight[36][98],
reservoir_weight[36][99],
reservoir_weight[36][100],
reservoir_weight[36][101],
reservoir_weight[36][102],
reservoir_weight[36][103],
reservoir_weight[36][104],
reservoir_weight[36][105],
reservoir_weight[36][106],
reservoir_weight[36][107],
reservoir_weight[36][108],
reservoir_weight[36][109],
reservoir_weight[36][110],
reservoir_weight[36][111],
reservoir_weight[36][112],
reservoir_weight[36][113],
reservoir_weight[36][114],
reservoir_weight[36][115],
reservoir_weight[36][116],
reservoir_weight[36][117],
reservoir_weight[36][118],
reservoir_weight[36][119],
reservoir_weight[36][120],
reservoir_weight[36][121],
reservoir_weight[36][122],
reservoir_weight[36][123],
reservoir_weight[36][124],
reservoir_weight[36][125],
reservoir_weight[36][126],
reservoir_weight[36][127],
reservoir_weight[36][128],
reservoir_weight[36][129],
reservoir_weight[36][130],
reservoir_weight[36][131],
reservoir_weight[36][132],
reservoir_weight[36][133],
reservoir_weight[36][134],
reservoir_weight[36][135],
reservoir_weight[36][136],
reservoir_weight[36][137],
reservoir_weight[36][138],
reservoir_weight[36][139],
reservoir_weight[36][140],
reservoir_weight[36][141],
reservoir_weight[36][142],
reservoir_weight[36][143],
reservoir_weight[36][144],
reservoir_weight[36][145],
reservoir_weight[36][146],
reservoir_weight[36][147],
reservoir_weight[36][148],
reservoir_weight[36][149],
reservoir_weight[36][150],
reservoir_weight[36][151],
reservoir_weight[36][152],
reservoir_weight[36][153],
reservoir_weight[36][154],
reservoir_weight[36][155],
reservoir_weight[36][156],
reservoir_weight[36][157],
reservoir_weight[36][158],
reservoir_weight[36][159],
reservoir_weight[36][160],
reservoir_weight[36][161],
reservoir_weight[36][162],
reservoir_weight[36][163],
reservoir_weight[36][164],
reservoir_weight[36][165],
reservoir_weight[36][166],
reservoir_weight[36][167],
reservoir_weight[36][168],
reservoir_weight[36][169],
reservoir_weight[36][170],
reservoir_weight[36][171],
reservoir_weight[36][172],
reservoir_weight[36][173],
reservoir_weight[36][174],
reservoir_weight[36][175],
reservoir_weight[36][176],
reservoir_weight[36][177],
reservoir_weight[36][178],
reservoir_weight[36][179],
reservoir_weight[36][180],
reservoir_weight[36][181],
reservoir_weight[36][182],
reservoir_weight[36][183],
reservoir_weight[36][184],
reservoir_weight[36][185],
reservoir_weight[36][186],
reservoir_weight[36][187],
reservoir_weight[36][188],
reservoir_weight[36][189],
reservoir_weight[36][190],
reservoir_weight[36][191],
reservoir_weight[36][192],
reservoir_weight[36][193],
reservoir_weight[36][194],
reservoir_weight[36][195],
reservoir_weight[36][196],
reservoir_weight[36][197],
reservoir_weight[36][198],
reservoir_weight[36][199]
},
{reservoir_weight[37][0],
reservoir_weight[37][1],
reservoir_weight[37][2],
reservoir_weight[37][3],
reservoir_weight[37][4],
reservoir_weight[37][5],
reservoir_weight[37][6],
reservoir_weight[37][7],
reservoir_weight[37][8],
reservoir_weight[37][9],
reservoir_weight[37][10],
reservoir_weight[37][11],
reservoir_weight[37][12],
reservoir_weight[37][13],
reservoir_weight[37][14],
reservoir_weight[37][15],
reservoir_weight[37][16],
reservoir_weight[37][17],
reservoir_weight[37][18],
reservoir_weight[37][19],
reservoir_weight[37][20],
reservoir_weight[37][21],
reservoir_weight[37][22],
reservoir_weight[37][23],
reservoir_weight[37][24],
reservoir_weight[37][25],
reservoir_weight[37][26],
reservoir_weight[37][27],
reservoir_weight[37][28],
reservoir_weight[37][29],
reservoir_weight[37][30],
reservoir_weight[37][31],
reservoir_weight[37][32],
reservoir_weight[37][33],
reservoir_weight[37][34],
reservoir_weight[37][35],
reservoir_weight[37][36],
reservoir_weight[37][37],
reservoir_weight[37][38],
reservoir_weight[37][39],
reservoir_weight[37][40],
reservoir_weight[37][41],
reservoir_weight[37][42],
reservoir_weight[37][43],
reservoir_weight[37][44],
reservoir_weight[37][45],
reservoir_weight[37][46],
reservoir_weight[37][47],
reservoir_weight[37][48],
reservoir_weight[37][49],
reservoir_weight[37][50],
reservoir_weight[37][51],
reservoir_weight[37][52],
reservoir_weight[37][53],
reservoir_weight[37][54],
reservoir_weight[37][55],
reservoir_weight[37][56],
reservoir_weight[37][57],
reservoir_weight[37][58],
reservoir_weight[37][59],
reservoir_weight[37][60],
reservoir_weight[37][61],
reservoir_weight[37][62],
reservoir_weight[37][63],
reservoir_weight[37][64],
reservoir_weight[37][65],
reservoir_weight[37][66],
reservoir_weight[37][67],
reservoir_weight[37][68],
reservoir_weight[37][69],
reservoir_weight[37][70],
reservoir_weight[37][71],
reservoir_weight[37][72],
reservoir_weight[37][73],
reservoir_weight[37][74],
reservoir_weight[37][75],
reservoir_weight[37][76],
reservoir_weight[37][77],
reservoir_weight[37][78],
reservoir_weight[37][79],
reservoir_weight[37][80],
reservoir_weight[37][81],
reservoir_weight[37][82],
reservoir_weight[37][83],
reservoir_weight[37][84],
reservoir_weight[37][85],
reservoir_weight[37][86],
reservoir_weight[37][87],
reservoir_weight[37][88],
reservoir_weight[37][89],
reservoir_weight[37][90],
reservoir_weight[37][91],
reservoir_weight[37][92],
reservoir_weight[37][93],
reservoir_weight[37][94],
reservoir_weight[37][95],
reservoir_weight[37][96],
reservoir_weight[37][97],
reservoir_weight[37][98],
reservoir_weight[37][99],
reservoir_weight[37][100],
reservoir_weight[37][101],
reservoir_weight[37][102],
reservoir_weight[37][103],
reservoir_weight[37][104],
reservoir_weight[37][105],
reservoir_weight[37][106],
reservoir_weight[37][107],
reservoir_weight[37][108],
reservoir_weight[37][109],
reservoir_weight[37][110],
reservoir_weight[37][111],
reservoir_weight[37][112],
reservoir_weight[37][113],
reservoir_weight[37][114],
reservoir_weight[37][115],
reservoir_weight[37][116],
reservoir_weight[37][117],
reservoir_weight[37][118],
reservoir_weight[37][119],
reservoir_weight[37][120],
reservoir_weight[37][121],
reservoir_weight[37][122],
reservoir_weight[37][123],
reservoir_weight[37][124],
reservoir_weight[37][125],
reservoir_weight[37][126],
reservoir_weight[37][127],
reservoir_weight[37][128],
reservoir_weight[37][129],
reservoir_weight[37][130],
reservoir_weight[37][131],
reservoir_weight[37][132],
reservoir_weight[37][133],
reservoir_weight[37][134],
reservoir_weight[37][135],
reservoir_weight[37][136],
reservoir_weight[37][137],
reservoir_weight[37][138],
reservoir_weight[37][139],
reservoir_weight[37][140],
reservoir_weight[37][141],
reservoir_weight[37][142],
reservoir_weight[37][143],
reservoir_weight[37][144],
reservoir_weight[37][145],
reservoir_weight[37][146],
reservoir_weight[37][147],
reservoir_weight[37][148],
reservoir_weight[37][149],
reservoir_weight[37][150],
reservoir_weight[37][151],
reservoir_weight[37][152],
reservoir_weight[37][153],
reservoir_weight[37][154],
reservoir_weight[37][155],
reservoir_weight[37][156],
reservoir_weight[37][157],
reservoir_weight[37][158],
reservoir_weight[37][159],
reservoir_weight[37][160],
reservoir_weight[37][161],
reservoir_weight[37][162],
reservoir_weight[37][163],
reservoir_weight[37][164],
reservoir_weight[37][165],
reservoir_weight[37][166],
reservoir_weight[37][167],
reservoir_weight[37][168],
reservoir_weight[37][169],
reservoir_weight[37][170],
reservoir_weight[37][171],
reservoir_weight[37][172],
reservoir_weight[37][173],
reservoir_weight[37][174],
reservoir_weight[37][175],
reservoir_weight[37][176],
reservoir_weight[37][177],
reservoir_weight[37][178],
reservoir_weight[37][179],
reservoir_weight[37][180],
reservoir_weight[37][181],
reservoir_weight[37][182],
reservoir_weight[37][183],
reservoir_weight[37][184],
reservoir_weight[37][185],
reservoir_weight[37][186],
reservoir_weight[37][187],
reservoir_weight[37][188],
reservoir_weight[37][189],
reservoir_weight[37][190],
reservoir_weight[37][191],
reservoir_weight[37][192],
reservoir_weight[37][193],
reservoir_weight[37][194],
reservoir_weight[37][195],
reservoir_weight[37][196],
reservoir_weight[37][197],
reservoir_weight[37][198],
reservoir_weight[37][199]
},
{reservoir_weight[38][0],
reservoir_weight[38][1],
reservoir_weight[38][2],
reservoir_weight[38][3],
reservoir_weight[38][4],
reservoir_weight[38][5],
reservoir_weight[38][6],
reservoir_weight[38][7],
reservoir_weight[38][8],
reservoir_weight[38][9],
reservoir_weight[38][10],
reservoir_weight[38][11],
reservoir_weight[38][12],
reservoir_weight[38][13],
reservoir_weight[38][14],
reservoir_weight[38][15],
reservoir_weight[38][16],
reservoir_weight[38][17],
reservoir_weight[38][18],
reservoir_weight[38][19],
reservoir_weight[38][20],
reservoir_weight[38][21],
reservoir_weight[38][22],
reservoir_weight[38][23],
reservoir_weight[38][24],
reservoir_weight[38][25],
reservoir_weight[38][26],
reservoir_weight[38][27],
reservoir_weight[38][28],
reservoir_weight[38][29],
reservoir_weight[38][30],
reservoir_weight[38][31],
reservoir_weight[38][32],
reservoir_weight[38][33],
reservoir_weight[38][34],
reservoir_weight[38][35],
reservoir_weight[38][36],
reservoir_weight[38][37],
reservoir_weight[38][38],
reservoir_weight[38][39],
reservoir_weight[38][40],
reservoir_weight[38][41],
reservoir_weight[38][42],
reservoir_weight[38][43],
reservoir_weight[38][44],
reservoir_weight[38][45],
reservoir_weight[38][46],
reservoir_weight[38][47],
reservoir_weight[38][48],
reservoir_weight[38][49],
reservoir_weight[38][50],
reservoir_weight[38][51],
reservoir_weight[38][52],
reservoir_weight[38][53],
reservoir_weight[38][54],
reservoir_weight[38][55],
reservoir_weight[38][56],
reservoir_weight[38][57],
reservoir_weight[38][58],
reservoir_weight[38][59],
reservoir_weight[38][60],
reservoir_weight[38][61],
reservoir_weight[38][62],
reservoir_weight[38][63],
reservoir_weight[38][64],
reservoir_weight[38][65],
reservoir_weight[38][66],
reservoir_weight[38][67],
reservoir_weight[38][68],
reservoir_weight[38][69],
reservoir_weight[38][70],
reservoir_weight[38][71],
reservoir_weight[38][72],
reservoir_weight[38][73],
reservoir_weight[38][74],
reservoir_weight[38][75],
reservoir_weight[38][76],
reservoir_weight[38][77],
reservoir_weight[38][78],
reservoir_weight[38][79],
reservoir_weight[38][80],
reservoir_weight[38][81],
reservoir_weight[38][82],
reservoir_weight[38][83],
reservoir_weight[38][84],
reservoir_weight[38][85],
reservoir_weight[38][86],
reservoir_weight[38][87],
reservoir_weight[38][88],
reservoir_weight[38][89],
reservoir_weight[38][90],
reservoir_weight[38][91],
reservoir_weight[38][92],
reservoir_weight[38][93],
reservoir_weight[38][94],
reservoir_weight[38][95],
reservoir_weight[38][96],
reservoir_weight[38][97],
reservoir_weight[38][98],
reservoir_weight[38][99],
reservoir_weight[38][100],
reservoir_weight[38][101],
reservoir_weight[38][102],
reservoir_weight[38][103],
reservoir_weight[38][104],
reservoir_weight[38][105],
reservoir_weight[38][106],
reservoir_weight[38][107],
reservoir_weight[38][108],
reservoir_weight[38][109],
reservoir_weight[38][110],
reservoir_weight[38][111],
reservoir_weight[38][112],
reservoir_weight[38][113],
reservoir_weight[38][114],
reservoir_weight[38][115],
reservoir_weight[38][116],
reservoir_weight[38][117],
reservoir_weight[38][118],
reservoir_weight[38][119],
reservoir_weight[38][120],
reservoir_weight[38][121],
reservoir_weight[38][122],
reservoir_weight[38][123],
reservoir_weight[38][124],
reservoir_weight[38][125],
reservoir_weight[38][126],
reservoir_weight[38][127],
reservoir_weight[38][128],
reservoir_weight[38][129],
reservoir_weight[38][130],
reservoir_weight[38][131],
reservoir_weight[38][132],
reservoir_weight[38][133],
reservoir_weight[38][134],
reservoir_weight[38][135],
reservoir_weight[38][136],
reservoir_weight[38][137],
reservoir_weight[38][138],
reservoir_weight[38][139],
reservoir_weight[38][140],
reservoir_weight[38][141],
reservoir_weight[38][142],
reservoir_weight[38][143],
reservoir_weight[38][144],
reservoir_weight[38][145],
reservoir_weight[38][146],
reservoir_weight[38][147],
reservoir_weight[38][148],
reservoir_weight[38][149],
reservoir_weight[38][150],
reservoir_weight[38][151],
reservoir_weight[38][152],
reservoir_weight[38][153],
reservoir_weight[38][154],
reservoir_weight[38][155],
reservoir_weight[38][156],
reservoir_weight[38][157],
reservoir_weight[38][158],
reservoir_weight[38][159],
reservoir_weight[38][160],
reservoir_weight[38][161],
reservoir_weight[38][162],
reservoir_weight[38][163],
reservoir_weight[38][164],
reservoir_weight[38][165],
reservoir_weight[38][166],
reservoir_weight[38][167],
reservoir_weight[38][168],
reservoir_weight[38][169],
reservoir_weight[38][170],
reservoir_weight[38][171],
reservoir_weight[38][172],
reservoir_weight[38][173],
reservoir_weight[38][174],
reservoir_weight[38][175],
reservoir_weight[38][176],
reservoir_weight[38][177],
reservoir_weight[38][178],
reservoir_weight[38][179],
reservoir_weight[38][180],
reservoir_weight[38][181],
reservoir_weight[38][182],
reservoir_weight[38][183],
reservoir_weight[38][184],
reservoir_weight[38][185],
reservoir_weight[38][186],
reservoir_weight[38][187],
reservoir_weight[38][188],
reservoir_weight[38][189],
reservoir_weight[38][190],
reservoir_weight[38][191],
reservoir_weight[38][192],
reservoir_weight[38][193],
reservoir_weight[38][194],
reservoir_weight[38][195],
reservoir_weight[38][196],
reservoir_weight[38][197],
reservoir_weight[38][198],
reservoir_weight[38][199]
},
{reservoir_weight[39][0],
reservoir_weight[39][1],
reservoir_weight[39][2],
reservoir_weight[39][3],
reservoir_weight[39][4],
reservoir_weight[39][5],
reservoir_weight[39][6],
reservoir_weight[39][7],
reservoir_weight[39][8],
reservoir_weight[39][9],
reservoir_weight[39][10],
reservoir_weight[39][11],
reservoir_weight[39][12],
reservoir_weight[39][13],
reservoir_weight[39][14],
reservoir_weight[39][15],
reservoir_weight[39][16],
reservoir_weight[39][17],
reservoir_weight[39][18],
reservoir_weight[39][19],
reservoir_weight[39][20],
reservoir_weight[39][21],
reservoir_weight[39][22],
reservoir_weight[39][23],
reservoir_weight[39][24],
reservoir_weight[39][25],
reservoir_weight[39][26],
reservoir_weight[39][27],
reservoir_weight[39][28],
reservoir_weight[39][29],
reservoir_weight[39][30],
reservoir_weight[39][31],
reservoir_weight[39][32],
reservoir_weight[39][33],
reservoir_weight[39][34],
reservoir_weight[39][35],
reservoir_weight[39][36],
reservoir_weight[39][37],
reservoir_weight[39][38],
reservoir_weight[39][39],
reservoir_weight[39][40],
reservoir_weight[39][41],
reservoir_weight[39][42],
reservoir_weight[39][43],
reservoir_weight[39][44],
reservoir_weight[39][45],
reservoir_weight[39][46],
reservoir_weight[39][47],
reservoir_weight[39][48],
reservoir_weight[39][49],
reservoir_weight[39][50],
reservoir_weight[39][51],
reservoir_weight[39][52],
reservoir_weight[39][53],
reservoir_weight[39][54],
reservoir_weight[39][55],
reservoir_weight[39][56],
reservoir_weight[39][57],
reservoir_weight[39][58],
reservoir_weight[39][59],
reservoir_weight[39][60],
reservoir_weight[39][61],
reservoir_weight[39][62],
reservoir_weight[39][63],
reservoir_weight[39][64],
reservoir_weight[39][65],
reservoir_weight[39][66],
reservoir_weight[39][67],
reservoir_weight[39][68],
reservoir_weight[39][69],
reservoir_weight[39][70],
reservoir_weight[39][71],
reservoir_weight[39][72],
reservoir_weight[39][73],
reservoir_weight[39][74],
reservoir_weight[39][75],
reservoir_weight[39][76],
reservoir_weight[39][77],
reservoir_weight[39][78],
reservoir_weight[39][79],
reservoir_weight[39][80],
reservoir_weight[39][81],
reservoir_weight[39][82],
reservoir_weight[39][83],
reservoir_weight[39][84],
reservoir_weight[39][85],
reservoir_weight[39][86],
reservoir_weight[39][87],
reservoir_weight[39][88],
reservoir_weight[39][89],
reservoir_weight[39][90],
reservoir_weight[39][91],
reservoir_weight[39][92],
reservoir_weight[39][93],
reservoir_weight[39][94],
reservoir_weight[39][95],
reservoir_weight[39][96],
reservoir_weight[39][97],
reservoir_weight[39][98],
reservoir_weight[39][99],
reservoir_weight[39][100],
reservoir_weight[39][101],
reservoir_weight[39][102],
reservoir_weight[39][103],
reservoir_weight[39][104],
reservoir_weight[39][105],
reservoir_weight[39][106],
reservoir_weight[39][107],
reservoir_weight[39][108],
reservoir_weight[39][109],
reservoir_weight[39][110],
reservoir_weight[39][111],
reservoir_weight[39][112],
reservoir_weight[39][113],
reservoir_weight[39][114],
reservoir_weight[39][115],
reservoir_weight[39][116],
reservoir_weight[39][117],
reservoir_weight[39][118],
reservoir_weight[39][119],
reservoir_weight[39][120],
reservoir_weight[39][121],
reservoir_weight[39][122],
reservoir_weight[39][123],
reservoir_weight[39][124],
reservoir_weight[39][125],
reservoir_weight[39][126],
reservoir_weight[39][127],
reservoir_weight[39][128],
reservoir_weight[39][129],
reservoir_weight[39][130],
reservoir_weight[39][131],
reservoir_weight[39][132],
reservoir_weight[39][133],
reservoir_weight[39][134],
reservoir_weight[39][135],
reservoir_weight[39][136],
reservoir_weight[39][137],
reservoir_weight[39][138],
reservoir_weight[39][139],
reservoir_weight[39][140],
reservoir_weight[39][141],
reservoir_weight[39][142],
reservoir_weight[39][143],
reservoir_weight[39][144],
reservoir_weight[39][145],
reservoir_weight[39][146],
reservoir_weight[39][147],
reservoir_weight[39][148],
reservoir_weight[39][149],
reservoir_weight[39][150],
reservoir_weight[39][151],
reservoir_weight[39][152],
reservoir_weight[39][153],
reservoir_weight[39][154],
reservoir_weight[39][155],
reservoir_weight[39][156],
reservoir_weight[39][157],
reservoir_weight[39][158],
reservoir_weight[39][159],
reservoir_weight[39][160],
reservoir_weight[39][161],
reservoir_weight[39][162],
reservoir_weight[39][163],
reservoir_weight[39][164],
reservoir_weight[39][165],
reservoir_weight[39][166],
reservoir_weight[39][167],
reservoir_weight[39][168],
reservoir_weight[39][169],
reservoir_weight[39][170],
reservoir_weight[39][171],
reservoir_weight[39][172],
reservoir_weight[39][173],
reservoir_weight[39][174],
reservoir_weight[39][175],
reservoir_weight[39][176],
reservoir_weight[39][177],
reservoir_weight[39][178],
reservoir_weight[39][179],
reservoir_weight[39][180],
reservoir_weight[39][181],
reservoir_weight[39][182],
reservoir_weight[39][183],
reservoir_weight[39][184],
reservoir_weight[39][185],
reservoir_weight[39][186],
reservoir_weight[39][187],
reservoir_weight[39][188],
reservoir_weight[39][189],
reservoir_weight[39][190],
reservoir_weight[39][191],
reservoir_weight[39][192],
reservoir_weight[39][193],
reservoir_weight[39][194],
reservoir_weight[39][195],
reservoir_weight[39][196],
reservoir_weight[39][197],
reservoir_weight[39][198],
reservoir_weight[39][199]
},
{reservoir_weight[40][0],
reservoir_weight[40][1],
reservoir_weight[40][2],
reservoir_weight[40][3],
reservoir_weight[40][4],
reservoir_weight[40][5],
reservoir_weight[40][6],
reservoir_weight[40][7],
reservoir_weight[40][8],
reservoir_weight[40][9],
reservoir_weight[40][10],
reservoir_weight[40][11],
reservoir_weight[40][12],
reservoir_weight[40][13],
reservoir_weight[40][14],
reservoir_weight[40][15],
reservoir_weight[40][16],
reservoir_weight[40][17],
reservoir_weight[40][18],
reservoir_weight[40][19],
reservoir_weight[40][20],
reservoir_weight[40][21],
reservoir_weight[40][22],
reservoir_weight[40][23],
reservoir_weight[40][24],
reservoir_weight[40][25],
reservoir_weight[40][26],
reservoir_weight[40][27],
reservoir_weight[40][28],
reservoir_weight[40][29],
reservoir_weight[40][30],
reservoir_weight[40][31],
reservoir_weight[40][32],
reservoir_weight[40][33],
reservoir_weight[40][34],
reservoir_weight[40][35],
reservoir_weight[40][36],
reservoir_weight[40][37],
reservoir_weight[40][38],
reservoir_weight[40][39],
reservoir_weight[40][40],
reservoir_weight[40][41],
reservoir_weight[40][42],
reservoir_weight[40][43],
reservoir_weight[40][44],
reservoir_weight[40][45],
reservoir_weight[40][46],
reservoir_weight[40][47],
reservoir_weight[40][48],
reservoir_weight[40][49],
reservoir_weight[40][50],
reservoir_weight[40][51],
reservoir_weight[40][52],
reservoir_weight[40][53],
reservoir_weight[40][54],
reservoir_weight[40][55],
reservoir_weight[40][56],
reservoir_weight[40][57],
reservoir_weight[40][58],
reservoir_weight[40][59],
reservoir_weight[40][60],
reservoir_weight[40][61],
reservoir_weight[40][62],
reservoir_weight[40][63],
reservoir_weight[40][64],
reservoir_weight[40][65],
reservoir_weight[40][66],
reservoir_weight[40][67],
reservoir_weight[40][68],
reservoir_weight[40][69],
reservoir_weight[40][70],
reservoir_weight[40][71],
reservoir_weight[40][72],
reservoir_weight[40][73],
reservoir_weight[40][74],
reservoir_weight[40][75],
reservoir_weight[40][76],
reservoir_weight[40][77],
reservoir_weight[40][78],
reservoir_weight[40][79],
reservoir_weight[40][80],
reservoir_weight[40][81],
reservoir_weight[40][82],
reservoir_weight[40][83],
reservoir_weight[40][84],
reservoir_weight[40][85],
reservoir_weight[40][86],
reservoir_weight[40][87],
reservoir_weight[40][88],
reservoir_weight[40][89],
reservoir_weight[40][90],
reservoir_weight[40][91],
reservoir_weight[40][92],
reservoir_weight[40][93],
reservoir_weight[40][94],
reservoir_weight[40][95],
reservoir_weight[40][96],
reservoir_weight[40][97],
reservoir_weight[40][98],
reservoir_weight[40][99],
reservoir_weight[40][100],
reservoir_weight[40][101],
reservoir_weight[40][102],
reservoir_weight[40][103],
reservoir_weight[40][104],
reservoir_weight[40][105],
reservoir_weight[40][106],
reservoir_weight[40][107],
reservoir_weight[40][108],
reservoir_weight[40][109],
reservoir_weight[40][110],
reservoir_weight[40][111],
reservoir_weight[40][112],
reservoir_weight[40][113],
reservoir_weight[40][114],
reservoir_weight[40][115],
reservoir_weight[40][116],
reservoir_weight[40][117],
reservoir_weight[40][118],
reservoir_weight[40][119],
reservoir_weight[40][120],
reservoir_weight[40][121],
reservoir_weight[40][122],
reservoir_weight[40][123],
reservoir_weight[40][124],
reservoir_weight[40][125],
reservoir_weight[40][126],
reservoir_weight[40][127],
reservoir_weight[40][128],
reservoir_weight[40][129],
reservoir_weight[40][130],
reservoir_weight[40][131],
reservoir_weight[40][132],
reservoir_weight[40][133],
reservoir_weight[40][134],
reservoir_weight[40][135],
reservoir_weight[40][136],
reservoir_weight[40][137],
reservoir_weight[40][138],
reservoir_weight[40][139],
reservoir_weight[40][140],
reservoir_weight[40][141],
reservoir_weight[40][142],
reservoir_weight[40][143],
reservoir_weight[40][144],
reservoir_weight[40][145],
reservoir_weight[40][146],
reservoir_weight[40][147],
reservoir_weight[40][148],
reservoir_weight[40][149],
reservoir_weight[40][150],
reservoir_weight[40][151],
reservoir_weight[40][152],
reservoir_weight[40][153],
reservoir_weight[40][154],
reservoir_weight[40][155],
reservoir_weight[40][156],
reservoir_weight[40][157],
reservoir_weight[40][158],
reservoir_weight[40][159],
reservoir_weight[40][160],
reservoir_weight[40][161],
reservoir_weight[40][162],
reservoir_weight[40][163],
reservoir_weight[40][164],
reservoir_weight[40][165],
reservoir_weight[40][166],
reservoir_weight[40][167],
reservoir_weight[40][168],
reservoir_weight[40][169],
reservoir_weight[40][170],
reservoir_weight[40][171],
reservoir_weight[40][172],
reservoir_weight[40][173],
reservoir_weight[40][174],
reservoir_weight[40][175],
reservoir_weight[40][176],
reservoir_weight[40][177],
reservoir_weight[40][178],
reservoir_weight[40][179],
reservoir_weight[40][180],
reservoir_weight[40][181],
reservoir_weight[40][182],
reservoir_weight[40][183],
reservoir_weight[40][184],
reservoir_weight[40][185],
reservoir_weight[40][186],
reservoir_weight[40][187],
reservoir_weight[40][188],
reservoir_weight[40][189],
reservoir_weight[40][190],
reservoir_weight[40][191],
reservoir_weight[40][192],
reservoir_weight[40][193],
reservoir_weight[40][194],
reservoir_weight[40][195],
reservoir_weight[40][196],
reservoir_weight[40][197],
reservoir_weight[40][198],
reservoir_weight[40][199]
},
{reservoir_weight[41][0],
reservoir_weight[41][1],
reservoir_weight[41][2],
reservoir_weight[41][3],
reservoir_weight[41][4],
reservoir_weight[41][5],
reservoir_weight[41][6],
reservoir_weight[41][7],
reservoir_weight[41][8],
reservoir_weight[41][9],
reservoir_weight[41][10],
reservoir_weight[41][11],
reservoir_weight[41][12],
reservoir_weight[41][13],
reservoir_weight[41][14],
reservoir_weight[41][15],
reservoir_weight[41][16],
reservoir_weight[41][17],
reservoir_weight[41][18],
reservoir_weight[41][19],
reservoir_weight[41][20],
reservoir_weight[41][21],
reservoir_weight[41][22],
reservoir_weight[41][23],
reservoir_weight[41][24],
reservoir_weight[41][25],
reservoir_weight[41][26],
reservoir_weight[41][27],
reservoir_weight[41][28],
reservoir_weight[41][29],
reservoir_weight[41][30],
reservoir_weight[41][31],
reservoir_weight[41][32],
reservoir_weight[41][33],
reservoir_weight[41][34],
reservoir_weight[41][35],
reservoir_weight[41][36],
reservoir_weight[41][37],
reservoir_weight[41][38],
reservoir_weight[41][39],
reservoir_weight[41][40],
reservoir_weight[41][41],
reservoir_weight[41][42],
reservoir_weight[41][43],
reservoir_weight[41][44],
reservoir_weight[41][45],
reservoir_weight[41][46],
reservoir_weight[41][47],
reservoir_weight[41][48],
reservoir_weight[41][49],
reservoir_weight[41][50],
reservoir_weight[41][51],
reservoir_weight[41][52],
reservoir_weight[41][53],
reservoir_weight[41][54],
reservoir_weight[41][55],
reservoir_weight[41][56],
reservoir_weight[41][57],
reservoir_weight[41][58],
reservoir_weight[41][59],
reservoir_weight[41][60],
reservoir_weight[41][61],
reservoir_weight[41][62],
reservoir_weight[41][63],
reservoir_weight[41][64],
reservoir_weight[41][65],
reservoir_weight[41][66],
reservoir_weight[41][67],
reservoir_weight[41][68],
reservoir_weight[41][69],
reservoir_weight[41][70],
reservoir_weight[41][71],
reservoir_weight[41][72],
reservoir_weight[41][73],
reservoir_weight[41][74],
reservoir_weight[41][75],
reservoir_weight[41][76],
reservoir_weight[41][77],
reservoir_weight[41][78],
reservoir_weight[41][79],
reservoir_weight[41][80],
reservoir_weight[41][81],
reservoir_weight[41][82],
reservoir_weight[41][83],
reservoir_weight[41][84],
reservoir_weight[41][85],
reservoir_weight[41][86],
reservoir_weight[41][87],
reservoir_weight[41][88],
reservoir_weight[41][89],
reservoir_weight[41][90],
reservoir_weight[41][91],
reservoir_weight[41][92],
reservoir_weight[41][93],
reservoir_weight[41][94],
reservoir_weight[41][95],
reservoir_weight[41][96],
reservoir_weight[41][97],
reservoir_weight[41][98],
reservoir_weight[41][99],
reservoir_weight[41][100],
reservoir_weight[41][101],
reservoir_weight[41][102],
reservoir_weight[41][103],
reservoir_weight[41][104],
reservoir_weight[41][105],
reservoir_weight[41][106],
reservoir_weight[41][107],
reservoir_weight[41][108],
reservoir_weight[41][109],
reservoir_weight[41][110],
reservoir_weight[41][111],
reservoir_weight[41][112],
reservoir_weight[41][113],
reservoir_weight[41][114],
reservoir_weight[41][115],
reservoir_weight[41][116],
reservoir_weight[41][117],
reservoir_weight[41][118],
reservoir_weight[41][119],
reservoir_weight[41][120],
reservoir_weight[41][121],
reservoir_weight[41][122],
reservoir_weight[41][123],
reservoir_weight[41][124],
reservoir_weight[41][125],
reservoir_weight[41][126],
reservoir_weight[41][127],
reservoir_weight[41][128],
reservoir_weight[41][129],
reservoir_weight[41][130],
reservoir_weight[41][131],
reservoir_weight[41][132],
reservoir_weight[41][133],
reservoir_weight[41][134],
reservoir_weight[41][135],
reservoir_weight[41][136],
reservoir_weight[41][137],
reservoir_weight[41][138],
reservoir_weight[41][139],
reservoir_weight[41][140],
reservoir_weight[41][141],
reservoir_weight[41][142],
reservoir_weight[41][143],
reservoir_weight[41][144],
reservoir_weight[41][145],
reservoir_weight[41][146],
reservoir_weight[41][147],
reservoir_weight[41][148],
reservoir_weight[41][149],
reservoir_weight[41][150],
reservoir_weight[41][151],
reservoir_weight[41][152],
reservoir_weight[41][153],
reservoir_weight[41][154],
reservoir_weight[41][155],
reservoir_weight[41][156],
reservoir_weight[41][157],
reservoir_weight[41][158],
reservoir_weight[41][159],
reservoir_weight[41][160],
reservoir_weight[41][161],
reservoir_weight[41][162],
reservoir_weight[41][163],
reservoir_weight[41][164],
reservoir_weight[41][165],
reservoir_weight[41][166],
reservoir_weight[41][167],
reservoir_weight[41][168],
reservoir_weight[41][169],
reservoir_weight[41][170],
reservoir_weight[41][171],
reservoir_weight[41][172],
reservoir_weight[41][173],
reservoir_weight[41][174],
reservoir_weight[41][175],
reservoir_weight[41][176],
reservoir_weight[41][177],
reservoir_weight[41][178],
reservoir_weight[41][179],
reservoir_weight[41][180],
reservoir_weight[41][181],
reservoir_weight[41][182],
reservoir_weight[41][183],
reservoir_weight[41][184],
reservoir_weight[41][185],
reservoir_weight[41][186],
reservoir_weight[41][187],
reservoir_weight[41][188],
reservoir_weight[41][189],
reservoir_weight[41][190],
reservoir_weight[41][191],
reservoir_weight[41][192],
reservoir_weight[41][193],
reservoir_weight[41][194],
reservoir_weight[41][195],
reservoir_weight[41][196],
reservoir_weight[41][197],
reservoir_weight[41][198],
reservoir_weight[41][199]
},
{reservoir_weight[42][0],
reservoir_weight[42][1],
reservoir_weight[42][2],
reservoir_weight[42][3],
reservoir_weight[42][4],
reservoir_weight[42][5],
reservoir_weight[42][6],
reservoir_weight[42][7],
reservoir_weight[42][8],
reservoir_weight[42][9],
reservoir_weight[42][10],
reservoir_weight[42][11],
reservoir_weight[42][12],
reservoir_weight[42][13],
reservoir_weight[42][14],
reservoir_weight[42][15],
reservoir_weight[42][16],
reservoir_weight[42][17],
reservoir_weight[42][18],
reservoir_weight[42][19],
reservoir_weight[42][20],
reservoir_weight[42][21],
reservoir_weight[42][22],
reservoir_weight[42][23],
reservoir_weight[42][24],
reservoir_weight[42][25],
reservoir_weight[42][26],
reservoir_weight[42][27],
reservoir_weight[42][28],
reservoir_weight[42][29],
reservoir_weight[42][30],
reservoir_weight[42][31],
reservoir_weight[42][32],
reservoir_weight[42][33],
reservoir_weight[42][34],
reservoir_weight[42][35],
reservoir_weight[42][36],
reservoir_weight[42][37],
reservoir_weight[42][38],
reservoir_weight[42][39],
reservoir_weight[42][40],
reservoir_weight[42][41],
reservoir_weight[42][42],
reservoir_weight[42][43],
reservoir_weight[42][44],
reservoir_weight[42][45],
reservoir_weight[42][46],
reservoir_weight[42][47],
reservoir_weight[42][48],
reservoir_weight[42][49],
reservoir_weight[42][50],
reservoir_weight[42][51],
reservoir_weight[42][52],
reservoir_weight[42][53],
reservoir_weight[42][54],
reservoir_weight[42][55],
reservoir_weight[42][56],
reservoir_weight[42][57],
reservoir_weight[42][58],
reservoir_weight[42][59],
reservoir_weight[42][60],
reservoir_weight[42][61],
reservoir_weight[42][62],
reservoir_weight[42][63],
reservoir_weight[42][64],
reservoir_weight[42][65],
reservoir_weight[42][66],
reservoir_weight[42][67],
reservoir_weight[42][68],
reservoir_weight[42][69],
reservoir_weight[42][70],
reservoir_weight[42][71],
reservoir_weight[42][72],
reservoir_weight[42][73],
reservoir_weight[42][74],
reservoir_weight[42][75],
reservoir_weight[42][76],
reservoir_weight[42][77],
reservoir_weight[42][78],
reservoir_weight[42][79],
reservoir_weight[42][80],
reservoir_weight[42][81],
reservoir_weight[42][82],
reservoir_weight[42][83],
reservoir_weight[42][84],
reservoir_weight[42][85],
reservoir_weight[42][86],
reservoir_weight[42][87],
reservoir_weight[42][88],
reservoir_weight[42][89],
reservoir_weight[42][90],
reservoir_weight[42][91],
reservoir_weight[42][92],
reservoir_weight[42][93],
reservoir_weight[42][94],
reservoir_weight[42][95],
reservoir_weight[42][96],
reservoir_weight[42][97],
reservoir_weight[42][98],
reservoir_weight[42][99],
reservoir_weight[42][100],
reservoir_weight[42][101],
reservoir_weight[42][102],
reservoir_weight[42][103],
reservoir_weight[42][104],
reservoir_weight[42][105],
reservoir_weight[42][106],
reservoir_weight[42][107],
reservoir_weight[42][108],
reservoir_weight[42][109],
reservoir_weight[42][110],
reservoir_weight[42][111],
reservoir_weight[42][112],
reservoir_weight[42][113],
reservoir_weight[42][114],
reservoir_weight[42][115],
reservoir_weight[42][116],
reservoir_weight[42][117],
reservoir_weight[42][118],
reservoir_weight[42][119],
reservoir_weight[42][120],
reservoir_weight[42][121],
reservoir_weight[42][122],
reservoir_weight[42][123],
reservoir_weight[42][124],
reservoir_weight[42][125],
reservoir_weight[42][126],
reservoir_weight[42][127],
reservoir_weight[42][128],
reservoir_weight[42][129],
reservoir_weight[42][130],
reservoir_weight[42][131],
reservoir_weight[42][132],
reservoir_weight[42][133],
reservoir_weight[42][134],
reservoir_weight[42][135],
reservoir_weight[42][136],
reservoir_weight[42][137],
reservoir_weight[42][138],
reservoir_weight[42][139],
reservoir_weight[42][140],
reservoir_weight[42][141],
reservoir_weight[42][142],
reservoir_weight[42][143],
reservoir_weight[42][144],
reservoir_weight[42][145],
reservoir_weight[42][146],
reservoir_weight[42][147],
reservoir_weight[42][148],
reservoir_weight[42][149],
reservoir_weight[42][150],
reservoir_weight[42][151],
reservoir_weight[42][152],
reservoir_weight[42][153],
reservoir_weight[42][154],
reservoir_weight[42][155],
reservoir_weight[42][156],
reservoir_weight[42][157],
reservoir_weight[42][158],
reservoir_weight[42][159],
reservoir_weight[42][160],
reservoir_weight[42][161],
reservoir_weight[42][162],
reservoir_weight[42][163],
reservoir_weight[42][164],
reservoir_weight[42][165],
reservoir_weight[42][166],
reservoir_weight[42][167],
reservoir_weight[42][168],
reservoir_weight[42][169],
reservoir_weight[42][170],
reservoir_weight[42][171],
reservoir_weight[42][172],
reservoir_weight[42][173],
reservoir_weight[42][174],
reservoir_weight[42][175],
reservoir_weight[42][176],
reservoir_weight[42][177],
reservoir_weight[42][178],
reservoir_weight[42][179],
reservoir_weight[42][180],
reservoir_weight[42][181],
reservoir_weight[42][182],
reservoir_weight[42][183],
reservoir_weight[42][184],
reservoir_weight[42][185],
reservoir_weight[42][186],
reservoir_weight[42][187],
reservoir_weight[42][188],
reservoir_weight[42][189],
reservoir_weight[42][190],
reservoir_weight[42][191],
reservoir_weight[42][192],
reservoir_weight[42][193],
reservoir_weight[42][194],
reservoir_weight[42][195],
reservoir_weight[42][196],
reservoir_weight[42][197],
reservoir_weight[42][198],
reservoir_weight[42][199]
},
{reservoir_weight[43][0],
reservoir_weight[43][1],
reservoir_weight[43][2],
reservoir_weight[43][3],
reservoir_weight[43][4],
reservoir_weight[43][5],
reservoir_weight[43][6],
reservoir_weight[43][7],
reservoir_weight[43][8],
reservoir_weight[43][9],
reservoir_weight[43][10],
reservoir_weight[43][11],
reservoir_weight[43][12],
reservoir_weight[43][13],
reservoir_weight[43][14],
reservoir_weight[43][15],
reservoir_weight[43][16],
reservoir_weight[43][17],
reservoir_weight[43][18],
reservoir_weight[43][19],
reservoir_weight[43][20],
reservoir_weight[43][21],
reservoir_weight[43][22],
reservoir_weight[43][23],
reservoir_weight[43][24],
reservoir_weight[43][25],
reservoir_weight[43][26],
reservoir_weight[43][27],
reservoir_weight[43][28],
reservoir_weight[43][29],
reservoir_weight[43][30],
reservoir_weight[43][31],
reservoir_weight[43][32],
reservoir_weight[43][33],
reservoir_weight[43][34],
reservoir_weight[43][35],
reservoir_weight[43][36],
reservoir_weight[43][37],
reservoir_weight[43][38],
reservoir_weight[43][39],
reservoir_weight[43][40],
reservoir_weight[43][41],
reservoir_weight[43][42],
reservoir_weight[43][43],
reservoir_weight[43][44],
reservoir_weight[43][45],
reservoir_weight[43][46],
reservoir_weight[43][47],
reservoir_weight[43][48],
reservoir_weight[43][49],
reservoir_weight[43][50],
reservoir_weight[43][51],
reservoir_weight[43][52],
reservoir_weight[43][53],
reservoir_weight[43][54],
reservoir_weight[43][55],
reservoir_weight[43][56],
reservoir_weight[43][57],
reservoir_weight[43][58],
reservoir_weight[43][59],
reservoir_weight[43][60],
reservoir_weight[43][61],
reservoir_weight[43][62],
reservoir_weight[43][63],
reservoir_weight[43][64],
reservoir_weight[43][65],
reservoir_weight[43][66],
reservoir_weight[43][67],
reservoir_weight[43][68],
reservoir_weight[43][69],
reservoir_weight[43][70],
reservoir_weight[43][71],
reservoir_weight[43][72],
reservoir_weight[43][73],
reservoir_weight[43][74],
reservoir_weight[43][75],
reservoir_weight[43][76],
reservoir_weight[43][77],
reservoir_weight[43][78],
reservoir_weight[43][79],
reservoir_weight[43][80],
reservoir_weight[43][81],
reservoir_weight[43][82],
reservoir_weight[43][83],
reservoir_weight[43][84],
reservoir_weight[43][85],
reservoir_weight[43][86],
reservoir_weight[43][87],
reservoir_weight[43][88],
reservoir_weight[43][89],
reservoir_weight[43][90],
reservoir_weight[43][91],
reservoir_weight[43][92],
reservoir_weight[43][93],
reservoir_weight[43][94],
reservoir_weight[43][95],
reservoir_weight[43][96],
reservoir_weight[43][97],
reservoir_weight[43][98],
reservoir_weight[43][99],
reservoir_weight[43][100],
reservoir_weight[43][101],
reservoir_weight[43][102],
reservoir_weight[43][103],
reservoir_weight[43][104],
reservoir_weight[43][105],
reservoir_weight[43][106],
reservoir_weight[43][107],
reservoir_weight[43][108],
reservoir_weight[43][109],
reservoir_weight[43][110],
reservoir_weight[43][111],
reservoir_weight[43][112],
reservoir_weight[43][113],
reservoir_weight[43][114],
reservoir_weight[43][115],
reservoir_weight[43][116],
reservoir_weight[43][117],
reservoir_weight[43][118],
reservoir_weight[43][119],
reservoir_weight[43][120],
reservoir_weight[43][121],
reservoir_weight[43][122],
reservoir_weight[43][123],
reservoir_weight[43][124],
reservoir_weight[43][125],
reservoir_weight[43][126],
reservoir_weight[43][127],
reservoir_weight[43][128],
reservoir_weight[43][129],
reservoir_weight[43][130],
reservoir_weight[43][131],
reservoir_weight[43][132],
reservoir_weight[43][133],
reservoir_weight[43][134],
reservoir_weight[43][135],
reservoir_weight[43][136],
reservoir_weight[43][137],
reservoir_weight[43][138],
reservoir_weight[43][139],
reservoir_weight[43][140],
reservoir_weight[43][141],
reservoir_weight[43][142],
reservoir_weight[43][143],
reservoir_weight[43][144],
reservoir_weight[43][145],
reservoir_weight[43][146],
reservoir_weight[43][147],
reservoir_weight[43][148],
reservoir_weight[43][149],
reservoir_weight[43][150],
reservoir_weight[43][151],
reservoir_weight[43][152],
reservoir_weight[43][153],
reservoir_weight[43][154],
reservoir_weight[43][155],
reservoir_weight[43][156],
reservoir_weight[43][157],
reservoir_weight[43][158],
reservoir_weight[43][159],
reservoir_weight[43][160],
reservoir_weight[43][161],
reservoir_weight[43][162],
reservoir_weight[43][163],
reservoir_weight[43][164],
reservoir_weight[43][165],
reservoir_weight[43][166],
reservoir_weight[43][167],
reservoir_weight[43][168],
reservoir_weight[43][169],
reservoir_weight[43][170],
reservoir_weight[43][171],
reservoir_weight[43][172],
reservoir_weight[43][173],
reservoir_weight[43][174],
reservoir_weight[43][175],
reservoir_weight[43][176],
reservoir_weight[43][177],
reservoir_weight[43][178],
reservoir_weight[43][179],
reservoir_weight[43][180],
reservoir_weight[43][181],
reservoir_weight[43][182],
reservoir_weight[43][183],
reservoir_weight[43][184],
reservoir_weight[43][185],
reservoir_weight[43][186],
reservoir_weight[43][187],
reservoir_weight[43][188],
reservoir_weight[43][189],
reservoir_weight[43][190],
reservoir_weight[43][191],
reservoir_weight[43][192],
reservoir_weight[43][193],
reservoir_weight[43][194],
reservoir_weight[43][195],
reservoir_weight[43][196],
reservoir_weight[43][197],
reservoir_weight[43][198],
reservoir_weight[43][199]
},
{reservoir_weight[44][0],
reservoir_weight[44][1],
reservoir_weight[44][2],
reservoir_weight[44][3],
reservoir_weight[44][4],
reservoir_weight[44][5],
reservoir_weight[44][6],
reservoir_weight[44][7],
reservoir_weight[44][8],
reservoir_weight[44][9],
reservoir_weight[44][10],
reservoir_weight[44][11],
reservoir_weight[44][12],
reservoir_weight[44][13],
reservoir_weight[44][14],
reservoir_weight[44][15],
reservoir_weight[44][16],
reservoir_weight[44][17],
reservoir_weight[44][18],
reservoir_weight[44][19],
reservoir_weight[44][20],
reservoir_weight[44][21],
reservoir_weight[44][22],
reservoir_weight[44][23],
reservoir_weight[44][24],
reservoir_weight[44][25],
reservoir_weight[44][26],
reservoir_weight[44][27],
reservoir_weight[44][28],
reservoir_weight[44][29],
reservoir_weight[44][30],
reservoir_weight[44][31],
reservoir_weight[44][32],
reservoir_weight[44][33],
reservoir_weight[44][34],
reservoir_weight[44][35],
reservoir_weight[44][36],
reservoir_weight[44][37],
reservoir_weight[44][38],
reservoir_weight[44][39],
reservoir_weight[44][40],
reservoir_weight[44][41],
reservoir_weight[44][42],
reservoir_weight[44][43],
reservoir_weight[44][44],
reservoir_weight[44][45],
reservoir_weight[44][46],
reservoir_weight[44][47],
reservoir_weight[44][48],
reservoir_weight[44][49],
reservoir_weight[44][50],
reservoir_weight[44][51],
reservoir_weight[44][52],
reservoir_weight[44][53],
reservoir_weight[44][54],
reservoir_weight[44][55],
reservoir_weight[44][56],
reservoir_weight[44][57],
reservoir_weight[44][58],
reservoir_weight[44][59],
reservoir_weight[44][60],
reservoir_weight[44][61],
reservoir_weight[44][62],
reservoir_weight[44][63],
reservoir_weight[44][64],
reservoir_weight[44][65],
reservoir_weight[44][66],
reservoir_weight[44][67],
reservoir_weight[44][68],
reservoir_weight[44][69],
reservoir_weight[44][70],
reservoir_weight[44][71],
reservoir_weight[44][72],
reservoir_weight[44][73],
reservoir_weight[44][74],
reservoir_weight[44][75],
reservoir_weight[44][76],
reservoir_weight[44][77],
reservoir_weight[44][78],
reservoir_weight[44][79],
reservoir_weight[44][80],
reservoir_weight[44][81],
reservoir_weight[44][82],
reservoir_weight[44][83],
reservoir_weight[44][84],
reservoir_weight[44][85],
reservoir_weight[44][86],
reservoir_weight[44][87],
reservoir_weight[44][88],
reservoir_weight[44][89],
reservoir_weight[44][90],
reservoir_weight[44][91],
reservoir_weight[44][92],
reservoir_weight[44][93],
reservoir_weight[44][94],
reservoir_weight[44][95],
reservoir_weight[44][96],
reservoir_weight[44][97],
reservoir_weight[44][98],
reservoir_weight[44][99],
reservoir_weight[44][100],
reservoir_weight[44][101],
reservoir_weight[44][102],
reservoir_weight[44][103],
reservoir_weight[44][104],
reservoir_weight[44][105],
reservoir_weight[44][106],
reservoir_weight[44][107],
reservoir_weight[44][108],
reservoir_weight[44][109],
reservoir_weight[44][110],
reservoir_weight[44][111],
reservoir_weight[44][112],
reservoir_weight[44][113],
reservoir_weight[44][114],
reservoir_weight[44][115],
reservoir_weight[44][116],
reservoir_weight[44][117],
reservoir_weight[44][118],
reservoir_weight[44][119],
reservoir_weight[44][120],
reservoir_weight[44][121],
reservoir_weight[44][122],
reservoir_weight[44][123],
reservoir_weight[44][124],
reservoir_weight[44][125],
reservoir_weight[44][126],
reservoir_weight[44][127],
reservoir_weight[44][128],
reservoir_weight[44][129],
reservoir_weight[44][130],
reservoir_weight[44][131],
reservoir_weight[44][132],
reservoir_weight[44][133],
reservoir_weight[44][134],
reservoir_weight[44][135],
reservoir_weight[44][136],
reservoir_weight[44][137],
reservoir_weight[44][138],
reservoir_weight[44][139],
reservoir_weight[44][140],
reservoir_weight[44][141],
reservoir_weight[44][142],
reservoir_weight[44][143],
reservoir_weight[44][144],
reservoir_weight[44][145],
reservoir_weight[44][146],
reservoir_weight[44][147],
reservoir_weight[44][148],
reservoir_weight[44][149],
reservoir_weight[44][150],
reservoir_weight[44][151],
reservoir_weight[44][152],
reservoir_weight[44][153],
reservoir_weight[44][154],
reservoir_weight[44][155],
reservoir_weight[44][156],
reservoir_weight[44][157],
reservoir_weight[44][158],
reservoir_weight[44][159],
reservoir_weight[44][160],
reservoir_weight[44][161],
reservoir_weight[44][162],
reservoir_weight[44][163],
reservoir_weight[44][164],
reservoir_weight[44][165],
reservoir_weight[44][166],
reservoir_weight[44][167],
reservoir_weight[44][168],
reservoir_weight[44][169],
reservoir_weight[44][170],
reservoir_weight[44][171],
reservoir_weight[44][172],
reservoir_weight[44][173],
reservoir_weight[44][174],
reservoir_weight[44][175],
reservoir_weight[44][176],
reservoir_weight[44][177],
reservoir_weight[44][178],
reservoir_weight[44][179],
reservoir_weight[44][180],
reservoir_weight[44][181],
reservoir_weight[44][182],
reservoir_weight[44][183],
reservoir_weight[44][184],
reservoir_weight[44][185],
reservoir_weight[44][186],
reservoir_weight[44][187],
reservoir_weight[44][188],
reservoir_weight[44][189],
reservoir_weight[44][190],
reservoir_weight[44][191],
reservoir_weight[44][192],
reservoir_weight[44][193],
reservoir_weight[44][194],
reservoir_weight[44][195],
reservoir_weight[44][196],
reservoir_weight[44][197],
reservoir_weight[44][198],
reservoir_weight[44][199]
},
{reservoir_weight[45][0],
reservoir_weight[45][1],
reservoir_weight[45][2],
reservoir_weight[45][3],
reservoir_weight[45][4],
reservoir_weight[45][5],
reservoir_weight[45][6],
reservoir_weight[45][7],
reservoir_weight[45][8],
reservoir_weight[45][9],
reservoir_weight[45][10],
reservoir_weight[45][11],
reservoir_weight[45][12],
reservoir_weight[45][13],
reservoir_weight[45][14],
reservoir_weight[45][15],
reservoir_weight[45][16],
reservoir_weight[45][17],
reservoir_weight[45][18],
reservoir_weight[45][19],
reservoir_weight[45][20],
reservoir_weight[45][21],
reservoir_weight[45][22],
reservoir_weight[45][23],
reservoir_weight[45][24],
reservoir_weight[45][25],
reservoir_weight[45][26],
reservoir_weight[45][27],
reservoir_weight[45][28],
reservoir_weight[45][29],
reservoir_weight[45][30],
reservoir_weight[45][31],
reservoir_weight[45][32],
reservoir_weight[45][33],
reservoir_weight[45][34],
reservoir_weight[45][35],
reservoir_weight[45][36],
reservoir_weight[45][37],
reservoir_weight[45][38],
reservoir_weight[45][39],
reservoir_weight[45][40],
reservoir_weight[45][41],
reservoir_weight[45][42],
reservoir_weight[45][43],
reservoir_weight[45][44],
reservoir_weight[45][45],
reservoir_weight[45][46],
reservoir_weight[45][47],
reservoir_weight[45][48],
reservoir_weight[45][49],
reservoir_weight[45][50],
reservoir_weight[45][51],
reservoir_weight[45][52],
reservoir_weight[45][53],
reservoir_weight[45][54],
reservoir_weight[45][55],
reservoir_weight[45][56],
reservoir_weight[45][57],
reservoir_weight[45][58],
reservoir_weight[45][59],
reservoir_weight[45][60],
reservoir_weight[45][61],
reservoir_weight[45][62],
reservoir_weight[45][63],
reservoir_weight[45][64],
reservoir_weight[45][65],
reservoir_weight[45][66],
reservoir_weight[45][67],
reservoir_weight[45][68],
reservoir_weight[45][69],
reservoir_weight[45][70],
reservoir_weight[45][71],
reservoir_weight[45][72],
reservoir_weight[45][73],
reservoir_weight[45][74],
reservoir_weight[45][75],
reservoir_weight[45][76],
reservoir_weight[45][77],
reservoir_weight[45][78],
reservoir_weight[45][79],
reservoir_weight[45][80],
reservoir_weight[45][81],
reservoir_weight[45][82],
reservoir_weight[45][83],
reservoir_weight[45][84],
reservoir_weight[45][85],
reservoir_weight[45][86],
reservoir_weight[45][87],
reservoir_weight[45][88],
reservoir_weight[45][89],
reservoir_weight[45][90],
reservoir_weight[45][91],
reservoir_weight[45][92],
reservoir_weight[45][93],
reservoir_weight[45][94],
reservoir_weight[45][95],
reservoir_weight[45][96],
reservoir_weight[45][97],
reservoir_weight[45][98],
reservoir_weight[45][99],
reservoir_weight[45][100],
reservoir_weight[45][101],
reservoir_weight[45][102],
reservoir_weight[45][103],
reservoir_weight[45][104],
reservoir_weight[45][105],
reservoir_weight[45][106],
reservoir_weight[45][107],
reservoir_weight[45][108],
reservoir_weight[45][109],
reservoir_weight[45][110],
reservoir_weight[45][111],
reservoir_weight[45][112],
reservoir_weight[45][113],
reservoir_weight[45][114],
reservoir_weight[45][115],
reservoir_weight[45][116],
reservoir_weight[45][117],
reservoir_weight[45][118],
reservoir_weight[45][119],
reservoir_weight[45][120],
reservoir_weight[45][121],
reservoir_weight[45][122],
reservoir_weight[45][123],
reservoir_weight[45][124],
reservoir_weight[45][125],
reservoir_weight[45][126],
reservoir_weight[45][127],
reservoir_weight[45][128],
reservoir_weight[45][129],
reservoir_weight[45][130],
reservoir_weight[45][131],
reservoir_weight[45][132],
reservoir_weight[45][133],
reservoir_weight[45][134],
reservoir_weight[45][135],
reservoir_weight[45][136],
reservoir_weight[45][137],
reservoir_weight[45][138],
reservoir_weight[45][139],
reservoir_weight[45][140],
reservoir_weight[45][141],
reservoir_weight[45][142],
reservoir_weight[45][143],
reservoir_weight[45][144],
reservoir_weight[45][145],
reservoir_weight[45][146],
reservoir_weight[45][147],
reservoir_weight[45][148],
reservoir_weight[45][149],
reservoir_weight[45][150],
reservoir_weight[45][151],
reservoir_weight[45][152],
reservoir_weight[45][153],
reservoir_weight[45][154],
reservoir_weight[45][155],
reservoir_weight[45][156],
reservoir_weight[45][157],
reservoir_weight[45][158],
reservoir_weight[45][159],
reservoir_weight[45][160],
reservoir_weight[45][161],
reservoir_weight[45][162],
reservoir_weight[45][163],
reservoir_weight[45][164],
reservoir_weight[45][165],
reservoir_weight[45][166],
reservoir_weight[45][167],
reservoir_weight[45][168],
reservoir_weight[45][169],
reservoir_weight[45][170],
reservoir_weight[45][171],
reservoir_weight[45][172],
reservoir_weight[45][173],
reservoir_weight[45][174],
reservoir_weight[45][175],
reservoir_weight[45][176],
reservoir_weight[45][177],
reservoir_weight[45][178],
reservoir_weight[45][179],
reservoir_weight[45][180],
reservoir_weight[45][181],
reservoir_weight[45][182],
reservoir_weight[45][183],
reservoir_weight[45][184],
reservoir_weight[45][185],
reservoir_weight[45][186],
reservoir_weight[45][187],
reservoir_weight[45][188],
reservoir_weight[45][189],
reservoir_weight[45][190],
reservoir_weight[45][191],
reservoir_weight[45][192],
reservoir_weight[45][193],
reservoir_weight[45][194],
reservoir_weight[45][195],
reservoir_weight[45][196],
reservoir_weight[45][197],
reservoir_weight[45][198],
reservoir_weight[45][199]
},
{reservoir_weight[46][0],
reservoir_weight[46][1],
reservoir_weight[46][2],
reservoir_weight[46][3],
reservoir_weight[46][4],
reservoir_weight[46][5],
reservoir_weight[46][6],
reservoir_weight[46][7],
reservoir_weight[46][8],
reservoir_weight[46][9],
reservoir_weight[46][10],
reservoir_weight[46][11],
reservoir_weight[46][12],
reservoir_weight[46][13],
reservoir_weight[46][14],
reservoir_weight[46][15],
reservoir_weight[46][16],
reservoir_weight[46][17],
reservoir_weight[46][18],
reservoir_weight[46][19],
reservoir_weight[46][20],
reservoir_weight[46][21],
reservoir_weight[46][22],
reservoir_weight[46][23],
reservoir_weight[46][24],
reservoir_weight[46][25],
reservoir_weight[46][26],
reservoir_weight[46][27],
reservoir_weight[46][28],
reservoir_weight[46][29],
reservoir_weight[46][30],
reservoir_weight[46][31],
reservoir_weight[46][32],
reservoir_weight[46][33],
reservoir_weight[46][34],
reservoir_weight[46][35],
reservoir_weight[46][36],
reservoir_weight[46][37],
reservoir_weight[46][38],
reservoir_weight[46][39],
reservoir_weight[46][40],
reservoir_weight[46][41],
reservoir_weight[46][42],
reservoir_weight[46][43],
reservoir_weight[46][44],
reservoir_weight[46][45],
reservoir_weight[46][46],
reservoir_weight[46][47],
reservoir_weight[46][48],
reservoir_weight[46][49],
reservoir_weight[46][50],
reservoir_weight[46][51],
reservoir_weight[46][52],
reservoir_weight[46][53],
reservoir_weight[46][54],
reservoir_weight[46][55],
reservoir_weight[46][56],
reservoir_weight[46][57],
reservoir_weight[46][58],
reservoir_weight[46][59],
reservoir_weight[46][60],
reservoir_weight[46][61],
reservoir_weight[46][62],
reservoir_weight[46][63],
reservoir_weight[46][64],
reservoir_weight[46][65],
reservoir_weight[46][66],
reservoir_weight[46][67],
reservoir_weight[46][68],
reservoir_weight[46][69],
reservoir_weight[46][70],
reservoir_weight[46][71],
reservoir_weight[46][72],
reservoir_weight[46][73],
reservoir_weight[46][74],
reservoir_weight[46][75],
reservoir_weight[46][76],
reservoir_weight[46][77],
reservoir_weight[46][78],
reservoir_weight[46][79],
reservoir_weight[46][80],
reservoir_weight[46][81],
reservoir_weight[46][82],
reservoir_weight[46][83],
reservoir_weight[46][84],
reservoir_weight[46][85],
reservoir_weight[46][86],
reservoir_weight[46][87],
reservoir_weight[46][88],
reservoir_weight[46][89],
reservoir_weight[46][90],
reservoir_weight[46][91],
reservoir_weight[46][92],
reservoir_weight[46][93],
reservoir_weight[46][94],
reservoir_weight[46][95],
reservoir_weight[46][96],
reservoir_weight[46][97],
reservoir_weight[46][98],
reservoir_weight[46][99],
reservoir_weight[46][100],
reservoir_weight[46][101],
reservoir_weight[46][102],
reservoir_weight[46][103],
reservoir_weight[46][104],
reservoir_weight[46][105],
reservoir_weight[46][106],
reservoir_weight[46][107],
reservoir_weight[46][108],
reservoir_weight[46][109],
reservoir_weight[46][110],
reservoir_weight[46][111],
reservoir_weight[46][112],
reservoir_weight[46][113],
reservoir_weight[46][114],
reservoir_weight[46][115],
reservoir_weight[46][116],
reservoir_weight[46][117],
reservoir_weight[46][118],
reservoir_weight[46][119],
reservoir_weight[46][120],
reservoir_weight[46][121],
reservoir_weight[46][122],
reservoir_weight[46][123],
reservoir_weight[46][124],
reservoir_weight[46][125],
reservoir_weight[46][126],
reservoir_weight[46][127],
reservoir_weight[46][128],
reservoir_weight[46][129],
reservoir_weight[46][130],
reservoir_weight[46][131],
reservoir_weight[46][132],
reservoir_weight[46][133],
reservoir_weight[46][134],
reservoir_weight[46][135],
reservoir_weight[46][136],
reservoir_weight[46][137],
reservoir_weight[46][138],
reservoir_weight[46][139],
reservoir_weight[46][140],
reservoir_weight[46][141],
reservoir_weight[46][142],
reservoir_weight[46][143],
reservoir_weight[46][144],
reservoir_weight[46][145],
reservoir_weight[46][146],
reservoir_weight[46][147],
reservoir_weight[46][148],
reservoir_weight[46][149],
reservoir_weight[46][150],
reservoir_weight[46][151],
reservoir_weight[46][152],
reservoir_weight[46][153],
reservoir_weight[46][154],
reservoir_weight[46][155],
reservoir_weight[46][156],
reservoir_weight[46][157],
reservoir_weight[46][158],
reservoir_weight[46][159],
reservoir_weight[46][160],
reservoir_weight[46][161],
reservoir_weight[46][162],
reservoir_weight[46][163],
reservoir_weight[46][164],
reservoir_weight[46][165],
reservoir_weight[46][166],
reservoir_weight[46][167],
reservoir_weight[46][168],
reservoir_weight[46][169],
reservoir_weight[46][170],
reservoir_weight[46][171],
reservoir_weight[46][172],
reservoir_weight[46][173],
reservoir_weight[46][174],
reservoir_weight[46][175],
reservoir_weight[46][176],
reservoir_weight[46][177],
reservoir_weight[46][178],
reservoir_weight[46][179],
reservoir_weight[46][180],
reservoir_weight[46][181],
reservoir_weight[46][182],
reservoir_weight[46][183],
reservoir_weight[46][184],
reservoir_weight[46][185],
reservoir_weight[46][186],
reservoir_weight[46][187],
reservoir_weight[46][188],
reservoir_weight[46][189],
reservoir_weight[46][190],
reservoir_weight[46][191],
reservoir_weight[46][192],
reservoir_weight[46][193],
reservoir_weight[46][194],
reservoir_weight[46][195],
reservoir_weight[46][196],
reservoir_weight[46][197],
reservoir_weight[46][198],
reservoir_weight[46][199]
},
{reservoir_weight[47][0],
reservoir_weight[47][1],
reservoir_weight[47][2],
reservoir_weight[47][3],
reservoir_weight[47][4],
reservoir_weight[47][5],
reservoir_weight[47][6],
reservoir_weight[47][7],
reservoir_weight[47][8],
reservoir_weight[47][9],
reservoir_weight[47][10],
reservoir_weight[47][11],
reservoir_weight[47][12],
reservoir_weight[47][13],
reservoir_weight[47][14],
reservoir_weight[47][15],
reservoir_weight[47][16],
reservoir_weight[47][17],
reservoir_weight[47][18],
reservoir_weight[47][19],
reservoir_weight[47][20],
reservoir_weight[47][21],
reservoir_weight[47][22],
reservoir_weight[47][23],
reservoir_weight[47][24],
reservoir_weight[47][25],
reservoir_weight[47][26],
reservoir_weight[47][27],
reservoir_weight[47][28],
reservoir_weight[47][29],
reservoir_weight[47][30],
reservoir_weight[47][31],
reservoir_weight[47][32],
reservoir_weight[47][33],
reservoir_weight[47][34],
reservoir_weight[47][35],
reservoir_weight[47][36],
reservoir_weight[47][37],
reservoir_weight[47][38],
reservoir_weight[47][39],
reservoir_weight[47][40],
reservoir_weight[47][41],
reservoir_weight[47][42],
reservoir_weight[47][43],
reservoir_weight[47][44],
reservoir_weight[47][45],
reservoir_weight[47][46],
reservoir_weight[47][47],
reservoir_weight[47][48],
reservoir_weight[47][49],
reservoir_weight[47][50],
reservoir_weight[47][51],
reservoir_weight[47][52],
reservoir_weight[47][53],
reservoir_weight[47][54],
reservoir_weight[47][55],
reservoir_weight[47][56],
reservoir_weight[47][57],
reservoir_weight[47][58],
reservoir_weight[47][59],
reservoir_weight[47][60],
reservoir_weight[47][61],
reservoir_weight[47][62],
reservoir_weight[47][63],
reservoir_weight[47][64],
reservoir_weight[47][65],
reservoir_weight[47][66],
reservoir_weight[47][67],
reservoir_weight[47][68],
reservoir_weight[47][69],
reservoir_weight[47][70],
reservoir_weight[47][71],
reservoir_weight[47][72],
reservoir_weight[47][73],
reservoir_weight[47][74],
reservoir_weight[47][75],
reservoir_weight[47][76],
reservoir_weight[47][77],
reservoir_weight[47][78],
reservoir_weight[47][79],
reservoir_weight[47][80],
reservoir_weight[47][81],
reservoir_weight[47][82],
reservoir_weight[47][83],
reservoir_weight[47][84],
reservoir_weight[47][85],
reservoir_weight[47][86],
reservoir_weight[47][87],
reservoir_weight[47][88],
reservoir_weight[47][89],
reservoir_weight[47][90],
reservoir_weight[47][91],
reservoir_weight[47][92],
reservoir_weight[47][93],
reservoir_weight[47][94],
reservoir_weight[47][95],
reservoir_weight[47][96],
reservoir_weight[47][97],
reservoir_weight[47][98],
reservoir_weight[47][99],
reservoir_weight[47][100],
reservoir_weight[47][101],
reservoir_weight[47][102],
reservoir_weight[47][103],
reservoir_weight[47][104],
reservoir_weight[47][105],
reservoir_weight[47][106],
reservoir_weight[47][107],
reservoir_weight[47][108],
reservoir_weight[47][109],
reservoir_weight[47][110],
reservoir_weight[47][111],
reservoir_weight[47][112],
reservoir_weight[47][113],
reservoir_weight[47][114],
reservoir_weight[47][115],
reservoir_weight[47][116],
reservoir_weight[47][117],
reservoir_weight[47][118],
reservoir_weight[47][119],
reservoir_weight[47][120],
reservoir_weight[47][121],
reservoir_weight[47][122],
reservoir_weight[47][123],
reservoir_weight[47][124],
reservoir_weight[47][125],
reservoir_weight[47][126],
reservoir_weight[47][127],
reservoir_weight[47][128],
reservoir_weight[47][129],
reservoir_weight[47][130],
reservoir_weight[47][131],
reservoir_weight[47][132],
reservoir_weight[47][133],
reservoir_weight[47][134],
reservoir_weight[47][135],
reservoir_weight[47][136],
reservoir_weight[47][137],
reservoir_weight[47][138],
reservoir_weight[47][139],
reservoir_weight[47][140],
reservoir_weight[47][141],
reservoir_weight[47][142],
reservoir_weight[47][143],
reservoir_weight[47][144],
reservoir_weight[47][145],
reservoir_weight[47][146],
reservoir_weight[47][147],
reservoir_weight[47][148],
reservoir_weight[47][149],
reservoir_weight[47][150],
reservoir_weight[47][151],
reservoir_weight[47][152],
reservoir_weight[47][153],
reservoir_weight[47][154],
reservoir_weight[47][155],
reservoir_weight[47][156],
reservoir_weight[47][157],
reservoir_weight[47][158],
reservoir_weight[47][159],
reservoir_weight[47][160],
reservoir_weight[47][161],
reservoir_weight[47][162],
reservoir_weight[47][163],
reservoir_weight[47][164],
reservoir_weight[47][165],
reservoir_weight[47][166],
reservoir_weight[47][167],
reservoir_weight[47][168],
reservoir_weight[47][169],
reservoir_weight[47][170],
reservoir_weight[47][171],
reservoir_weight[47][172],
reservoir_weight[47][173],
reservoir_weight[47][174],
reservoir_weight[47][175],
reservoir_weight[47][176],
reservoir_weight[47][177],
reservoir_weight[47][178],
reservoir_weight[47][179],
reservoir_weight[47][180],
reservoir_weight[47][181],
reservoir_weight[47][182],
reservoir_weight[47][183],
reservoir_weight[47][184],
reservoir_weight[47][185],
reservoir_weight[47][186],
reservoir_weight[47][187],
reservoir_weight[47][188],
reservoir_weight[47][189],
reservoir_weight[47][190],
reservoir_weight[47][191],
reservoir_weight[47][192],
reservoir_weight[47][193],
reservoir_weight[47][194],
reservoir_weight[47][195],
reservoir_weight[47][196],
reservoir_weight[47][197],
reservoir_weight[47][198],
reservoir_weight[47][199]
},
{reservoir_weight[48][0],
reservoir_weight[48][1],
reservoir_weight[48][2],
reservoir_weight[48][3],
reservoir_weight[48][4],
reservoir_weight[48][5],
reservoir_weight[48][6],
reservoir_weight[48][7],
reservoir_weight[48][8],
reservoir_weight[48][9],
reservoir_weight[48][10],
reservoir_weight[48][11],
reservoir_weight[48][12],
reservoir_weight[48][13],
reservoir_weight[48][14],
reservoir_weight[48][15],
reservoir_weight[48][16],
reservoir_weight[48][17],
reservoir_weight[48][18],
reservoir_weight[48][19],
reservoir_weight[48][20],
reservoir_weight[48][21],
reservoir_weight[48][22],
reservoir_weight[48][23],
reservoir_weight[48][24],
reservoir_weight[48][25],
reservoir_weight[48][26],
reservoir_weight[48][27],
reservoir_weight[48][28],
reservoir_weight[48][29],
reservoir_weight[48][30],
reservoir_weight[48][31],
reservoir_weight[48][32],
reservoir_weight[48][33],
reservoir_weight[48][34],
reservoir_weight[48][35],
reservoir_weight[48][36],
reservoir_weight[48][37],
reservoir_weight[48][38],
reservoir_weight[48][39],
reservoir_weight[48][40],
reservoir_weight[48][41],
reservoir_weight[48][42],
reservoir_weight[48][43],
reservoir_weight[48][44],
reservoir_weight[48][45],
reservoir_weight[48][46],
reservoir_weight[48][47],
reservoir_weight[48][48],
reservoir_weight[48][49],
reservoir_weight[48][50],
reservoir_weight[48][51],
reservoir_weight[48][52],
reservoir_weight[48][53],
reservoir_weight[48][54],
reservoir_weight[48][55],
reservoir_weight[48][56],
reservoir_weight[48][57],
reservoir_weight[48][58],
reservoir_weight[48][59],
reservoir_weight[48][60],
reservoir_weight[48][61],
reservoir_weight[48][62],
reservoir_weight[48][63],
reservoir_weight[48][64],
reservoir_weight[48][65],
reservoir_weight[48][66],
reservoir_weight[48][67],
reservoir_weight[48][68],
reservoir_weight[48][69],
reservoir_weight[48][70],
reservoir_weight[48][71],
reservoir_weight[48][72],
reservoir_weight[48][73],
reservoir_weight[48][74],
reservoir_weight[48][75],
reservoir_weight[48][76],
reservoir_weight[48][77],
reservoir_weight[48][78],
reservoir_weight[48][79],
reservoir_weight[48][80],
reservoir_weight[48][81],
reservoir_weight[48][82],
reservoir_weight[48][83],
reservoir_weight[48][84],
reservoir_weight[48][85],
reservoir_weight[48][86],
reservoir_weight[48][87],
reservoir_weight[48][88],
reservoir_weight[48][89],
reservoir_weight[48][90],
reservoir_weight[48][91],
reservoir_weight[48][92],
reservoir_weight[48][93],
reservoir_weight[48][94],
reservoir_weight[48][95],
reservoir_weight[48][96],
reservoir_weight[48][97],
reservoir_weight[48][98],
reservoir_weight[48][99],
reservoir_weight[48][100],
reservoir_weight[48][101],
reservoir_weight[48][102],
reservoir_weight[48][103],
reservoir_weight[48][104],
reservoir_weight[48][105],
reservoir_weight[48][106],
reservoir_weight[48][107],
reservoir_weight[48][108],
reservoir_weight[48][109],
reservoir_weight[48][110],
reservoir_weight[48][111],
reservoir_weight[48][112],
reservoir_weight[48][113],
reservoir_weight[48][114],
reservoir_weight[48][115],
reservoir_weight[48][116],
reservoir_weight[48][117],
reservoir_weight[48][118],
reservoir_weight[48][119],
reservoir_weight[48][120],
reservoir_weight[48][121],
reservoir_weight[48][122],
reservoir_weight[48][123],
reservoir_weight[48][124],
reservoir_weight[48][125],
reservoir_weight[48][126],
reservoir_weight[48][127],
reservoir_weight[48][128],
reservoir_weight[48][129],
reservoir_weight[48][130],
reservoir_weight[48][131],
reservoir_weight[48][132],
reservoir_weight[48][133],
reservoir_weight[48][134],
reservoir_weight[48][135],
reservoir_weight[48][136],
reservoir_weight[48][137],
reservoir_weight[48][138],
reservoir_weight[48][139],
reservoir_weight[48][140],
reservoir_weight[48][141],
reservoir_weight[48][142],
reservoir_weight[48][143],
reservoir_weight[48][144],
reservoir_weight[48][145],
reservoir_weight[48][146],
reservoir_weight[48][147],
reservoir_weight[48][148],
reservoir_weight[48][149],
reservoir_weight[48][150],
reservoir_weight[48][151],
reservoir_weight[48][152],
reservoir_weight[48][153],
reservoir_weight[48][154],
reservoir_weight[48][155],
reservoir_weight[48][156],
reservoir_weight[48][157],
reservoir_weight[48][158],
reservoir_weight[48][159],
reservoir_weight[48][160],
reservoir_weight[48][161],
reservoir_weight[48][162],
reservoir_weight[48][163],
reservoir_weight[48][164],
reservoir_weight[48][165],
reservoir_weight[48][166],
reservoir_weight[48][167],
reservoir_weight[48][168],
reservoir_weight[48][169],
reservoir_weight[48][170],
reservoir_weight[48][171],
reservoir_weight[48][172],
reservoir_weight[48][173],
reservoir_weight[48][174],
reservoir_weight[48][175],
reservoir_weight[48][176],
reservoir_weight[48][177],
reservoir_weight[48][178],
reservoir_weight[48][179],
reservoir_weight[48][180],
reservoir_weight[48][181],
reservoir_weight[48][182],
reservoir_weight[48][183],
reservoir_weight[48][184],
reservoir_weight[48][185],
reservoir_weight[48][186],
reservoir_weight[48][187],
reservoir_weight[48][188],
reservoir_weight[48][189],
reservoir_weight[48][190],
reservoir_weight[48][191],
reservoir_weight[48][192],
reservoir_weight[48][193],
reservoir_weight[48][194],
reservoir_weight[48][195],
reservoir_weight[48][196],
reservoir_weight[48][197],
reservoir_weight[48][198],
reservoir_weight[48][199]
},
{reservoir_weight[49][0],
reservoir_weight[49][1],
reservoir_weight[49][2],
reservoir_weight[49][3],
reservoir_weight[49][4],
reservoir_weight[49][5],
reservoir_weight[49][6],
reservoir_weight[49][7],
reservoir_weight[49][8],
reservoir_weight[49][9],
reservoir_weight[49][10],
reservoir_weight[49][11],
reservoir_weight[49][12],
reservoir_weight[49][13],
reservoir_weight[49][14],
reservoir_weight[49][15],
reservoir_weight[49][16],
reservoir_weight[49][17],
reservoir_weight[49][18],
reservoir_weight[49][19],
reservoir_weight[49][20],
reservoir_weight[49][21],
reservoir_weight[49][22],
reservoir_weight[49][23],
reservoir_weight[49][24],
reservoir_weight[49][25],
reservoir_weight[49][26],
reservoir_weight[49][27],
reservoir_weight[49][28],
reservoir_weight[49][29],
reservoir_weight[49][30],
reservoir_weight[49][31],
reservoir_weight[49][32],
reservoir_weight[49][33],
reservoir_weight[49][34],
reservoir_weight[49][35],
reservoir_weight[49][36],
reservoir_weight[49][37],
reservoir_weight[49][38],
reservoir_weight[49][39],
reservoir_weight[49][40],
reservoir_weight[49][41],
reservoir_weight[49][42],
reservoir_weight[49][43],
reservoir_weight[49][44],
reservoir_weight[49][45],
reservoir_weight[49][46],
reservoir_weight[49][47],
reservoir_weight[49][48],
reservoir_weight[49][49],
reservoir_weight[49][50],
reservoir_weight[49][51],
reservoir_weight[49][52],
reservoir_weight[49][53],
reservoir_weight[49][54],
reservoir_weight[49][55],
reservoir_weight[49][56],
reservoir_weight[49][57],
reservoir_weight[49][58],
reservoir_weight[49][59],
reservoir_weight[49][60],
reservoir_weight[49][61],
reservoir_weight[49][62],
reservoir_weight[49][63],
reservoir_weight[49][64],
reservoir_weight[49][65],
reservoir_weight[49][66],
reservoir_weight[49][67],
reservoir_weight[49][68],
reservoir_weight[49][69],
reservoir_weight[49][70],
reservoir_weight[49][71],
reservoir_weight[49][72],
reservoir_weight[49][73],
reservoir_weight[49][74],
reservoir_weight[49][75],
reservoir_weight[49][76],
reservoir_weight[49][77],
reservoir_weight[49][78],
reservoir_weight[49][79],
reservoir_weight[49][80],
reservoir_weight[49][81],
reservoir_weight[49][82],
reservoir_weight[49][83],
reservoir_weight[49][84],
reservoir_weight[49][85],
reservoir_weight[49][86],
reservoir_weight[49][87],
reservoir_weight[49][88],
reservoir_weight[49][89],
reservoir_weight[49][90],
reservoir_weight[49][91],
reservoir_weight[49][92],
reservoir_weight[49][93],
reservoir_weight[49][94],
reservoir_weight[49][95],
reservoir_weight[49][96],
reservoir_weight[49][97],
reservoir_weight[49][98],
reservoir_weight[49][99],
reservoir_weight[49][100],
reservoir_weight[49][101],
reservoir_weight[49][102],
reservoir_weight[49][103],
reservoir_weight[49][104],
reservoir_weight[49][105],
reservoir_weight[49][106],
reservoir_weight[49][107],
reservoir_weight[49][108],
reservoir_weight[49][109],
reservoir_weight[49][110],
reservoir_weight[49][111],
reservoir_weight[49][112],
reservoir_weight[49][113],
reservoir_weight[49][114],
reservoir_weight[49][115],
reservoir_weight[49][116],
reservoir_weight[49][117],
reservoir_weight[49][118],
reservoir_weight[49][119],
reservoir_weight[49][120],
reservoir_weight[49][121],
reservoir_weight[49][122],
reservoir_weight[49][123],
reservoir_weight[49][124],
reservoir_weight[49][125],
reservoir_weight[49][126],
reservoir_weight[49][127],
reservoir_weight[49][128],
reservoir_weight[49][129],
reservoir_weight[49][130],
reservoir_weight[49][131],
reservoir_weight[49][132],
reservoir_weight[49][133],
reservoir_weight[49][134],
reservoir_weight[49][135],
reservoir_weight[49][136],
reservoir_weight[49][137],
reservoir_weight[49][138],
reservoir_weight[49][139],
reservoir_weight[49][140],
reservoir_weight[49][141],
reservoir_weight[49][142],
reservoir_weight[49][143],
reservoir_weight[49][144],
reservoir_weight[49][145],
reservoir_weight[49][146],
reservoir_weight[49][147],
reservoir_weight[49][148],
reservoir_weight[49][149],
reservoir_weight[49][150],
reservoir_weight[49][151],
reservoir_weight[49][152],
reservoir_weight[49][153],
reservoir_weight[49][154],
reservoir_weight[49][155],
reservoir_weight[49][156],
reservoir_weight[49][157],
reservoir_weight[49][158],
reservoir_weight[49][159],
reservoir_weight[49][160],
reservoir_weight[49][161],
reservoir_weight[49][162],
reservoir_weight[49][163],
reservoir_weight[49][164],
reservoir_weight[49][165],
reservoir_weight[49][166],
reservoir_weight[49][167],
reservoir_weight[49][168],
reservoir_weight[49][169],
reservoir_weight[49][170],
reservoir_weight[49][171],
reservoir_weight[49][172],
reservoir_weight[49][173],
reservoir_weight[49][174],
reservoir_weight[49][175],
reservoir_weight[49][176],
reservoir_weight[49][177],
reservoir_weight[49][178],
reservoir_weight[49][179],
reservoir_weight[49][180],
reservoir_weight[49][181],
reservoir_weight[49][182],
reservoir_weight[49][183],
reservoir_weight[49][184],
reservoir_weight[49][185],
reservoir_weight[49][186],
reservoir_weight[49][187],
reservoir_weight[49][188],
reservoir_weight[49][189],
reservoir_weight[49][190],
reservoir_weight[49][191],
reservoir_weight[49][192],
reservoir_weight[49][193],
reservoir_weight[49][194],
reservoir_weight[49][195],
reservoir_weight[49][196],
reservoir_weight[49][197],
reservoir_weight[49][198],
reservoir_weight[49][199]
},
{reservoir_weight[50][0],
reservoir_weight[50][1],
reservoir_weight[50][2],
reservoir_weight[50][3],
reservoir_weight[50][4],
reservoir_weight[50][5],
reservoir_weight[50][6],
reservoir_weight[50][7],
reservoir_weight[50][8],
reservoir_weight[50][9],
reservoir_weight[50][10],
reservoir_weight[50][11],
reservoir_weight[50][12],
reservoir_weight[50][13],
reservoir_weight[50][14],
reservoir_weight[50][15],
reservoir_weight[50][16],
reservoir_weight[50][17],
reservoir_weight[50][18],
reservoir_weight[50][19],
reservoir_weight[50][20],
reservoir_weight[50][21],
reservoir_weight[50][22],
reservoir_weight[50][23],
reservoir_weight[50][24],
reservoir_weight[50][25],
reservoir_weight[50][26],
reservoir_weight[50][27],
reservoir_weight[50][28],
reservoir_weight[50][29],
reservoir_weight[50][30],
reservoir_weight[50][31],
reservoir_weight[50][32],
reservoir_weight[50][33],
reservoir_weight[50][34],
reservoir_weight[50][35],
reservoir_weight[50][36],
reservoir_weight[50][37],
reservoir_weight[50][38],
reservoir_weight[50][39],
reservoir_weight[50][40],
reservoir_weight[50][41],
reservoir_weight[50][42],
reservoir_weight[50][43],
reservoir_weight[50][44],
reservoir_weight[50][45],
reservoir_weight[50][46],
reservoir_weight[50][47],
reservoir_weight[50][48],
reservoir_weight[50][49],
reservoir_weight[50][50],
reservoir_weight[50][51],
reservoir_weight[50][52],
reservoir_weight[50][53],
reservoir_weight[50][54],
reservoir_weight[50][55],
reservoir_weight[50][56],
reservoir_weight[50][57],
reservoir_weight[50][58],
reservoir_weight[50][59],
reservoir_weight[50][60],
reservoir_weight[50][61],
reservoir_weight[50][62],
reservoir_weight[50][63],
reservoir_weight[50][64],
reservoir_weight[50][65],
reservoir_weight[50][66],
reservoir_weight[50][67],
reservoir_weight[50][68],
reservoir_weight[50][69],
reservoir_weight[50][70],
reservoir_weight[50][71],
reservoir_weight[50][72],
reservoir_weight[50][73],
reservoir_weight[50][74],
reservoir_weight[50][75],
reservoir_weight[50][76],
reservoir_weight[50][77],
reservoir_weight[50][78],
reservoir_weight[50][79],
reservoir_weight[50][80],
reservoir_weight[50][81],
reservoir_weight[50][82],
reservoir_weight[50][83],
reservoir_weight[50][84],
reservoir_weight[50][85],
reservoir_weight[50][86],
reservoir_weight[50][87],
reservoir_weight[50][88],
reservoir_weight[50][89],
reservoir_weight[50][90],
reservoir_weight[50][91],
reservoir_weight[50][92],
reservoir_weight[50][93],
reservoir_weight[50][94],
reservoir_weight[50][95],
reservoir_weight[50][96],
reservoir_weight[50][97],
reservoir_weight[50][98],
reservoir_weight[50][99],
reservoir_weight[50][100],
reservoir_weight[50][101],
reservoir_weight[50][102],
reservoir_weight[50][103],
reservoir_weight[50][104],
reservoir_weight[50][105],
reservoir_weight[50][106],
reservoir_weight[50][107],
reservoir_weight[50][108],
reservoir_weight[50][109],
reservoir_weight[50][110],
reservoir_weight[50][111],
reservoir_weight[50][112],
reservoir_weight[50][113],
reservoir_weight[50][114],
reservoir_weight[50][115],
reservoir_weight[50][116],
reservoir_weight[50][117],
reservoir_weight[50][118],
reservoir_weight[50][119],
reservoir_weight[50][120],
reservoir_weight[50][121],
reservoir_weight[50][122],
reservoir_weight[50][123],
reservoir_weight[50][124],
reservoir_weight[50][125],
reservoir_weight[50][126],
reservoir_weight[50][127],
reservoir_weight[50][128],
reservoir_weight[50][129],
reservoir_weight[50][130],
reservoir_weight[50][131],
reservoir_weight[50][132],
reservoir_weight[50][133],
reservoir_weight[50][134],
reservoir_weight[50][135],
reservoir_weight[50][136],
reservoir_weight[50][137],
reservoir_weight[50][138],
reservoir_weight[50][139],
reservoir_weight[50][140],
reservoir_weight[50][141],
reservoir_weight[50][142],
reservoir_weight[50][143],
reservoir_weight[50][144],
reservoir_weight[50][145],
reservoir_weight[50][146],
reservoir_weight[50][147],
reservoir_weight[50][148],
reservoir_weight[50][149],
reservoir_weight[50][150],
reservoir_weight[50][151],
reservoir_weight[50][152],
reservoir_weight[50][153],
reservoir_weight[50][154],
reservoir_weight[50][155],
reservoir_weight[50][156],
reservoir_weight[50][157],
reservoir_weight[50][158],
reservoir_weight[50][159],
reservoir_weight[50][160],
reservoir_weight[50][161],
reservoir_weight[50][162],
reservoir_weight[50][163],
reservoir_weight[50][164],
reservoir_weight[50][165],
reservoir_weight[50][166],
reservoir_weight[50][167],
reservoir_weight[50][168],
reservoir_weight[50][169],
reservoir_weight[50][170],
reservoir_weight[50][171],
reservoir_weight[50][172],
reservoir_weight[50][173],
reservoir_weight[50][174],
reservoir_weight[50][175],
reservoir_weight[50][176],
reservoir_weight[50][177],
reservoir_weight[50][178],
reservoir_weight[50][179],
reservoir_weight[50][180],
reservoir_weight[50][181],
reservoir_weight[50][182],
reservoir_weight[50][183],
reservoir_weight[50][184],
reservoir_weight[50][185],
reservoir_weight[50][186],
reservoir_weight[50][187],
reservoir_weight[50][188],
reservoir_weight[50][189],
reservoir_weight[50][190],
reservoir_weight[50][191],
reservoir_weight[50][192],
reservoir_weight[50][193],
reservoir_weight[50][194],
reservoir_weight[50][195],
reservoir_weight[50][196],
reservoir_weight[50][197],
reservoir_weight[50][198],
reservoir_weight[50][199]
},
{reservoir_weight[51][0],
reservoir_weight[51][1],
reservoir_weight[51][2],
reservoir_weight[51][3],
reservoir_weight[51][4],
reservoir_weight[51][5],
reservoir_weight[51][6],
reservoir_weight[51][7],
reservoir_weight[51][8],
reservoir_weight[51][9],
reservoir_weight[51][10],
reservoir_weight[51][11],
reservoir_weight[51][12],
reservoir_weight[51][13],
reservoir_weight[51][14],
reservoir_weight[51][15],
reservoir_weight[51][16],
reservoir_weight[51][17],
reservoir_weight[51][18],
reservoir_weight[51][19],
reservoir_weight[51][20],
reservoir_weight[51][21],
reservoir_weight[51][22],
reservoir_weight[51][23],
reservoir_weight[51][24],
reservoir_weight[51][25],
reservoir_weight[51][26],
reservoir_weight[51][27],
reservoir_weight[51][28],
reservoir_weight[51][29],
reservoir_weight[51][30],
reservoir_weight[51][31],
reservoir_weight[51][32],
reservoir_weight[51][33],
reservoir_weight[51][34],
reservoir_weight[51][35],
reservoir_weight[51][36],
reservoir_weight[51][37],
reservoir_weight[51][38],
reservoir_weight[51][39],
reservoir_weight[51][40],
reservoir_weight[51][41],
reservoir_weight[51][42],
reservoir_weight[51][43],
reservoir_weight[51][44],
reservoir_weight[51][45],
reservoir_weight[51][46],
reservoir_weight[51][47],
reservoir_weight[51][48],
reservoir_weight[51][49],
reservoir_weight[51][50],
reservoir_weight[51][51],
reservoir_weight[51][52],
reservoir_weight[51][53],
reservoir_weight[51][54],
reservoir_weight[51][55],
reservoir_weight[51][56],
reservoir_weight[51][57],
reservoir_weight[51][58],
reservoir_weight[51][59],
reservoir_weight[51][60],
reservoir_weight[51][61],
reservoir_weight[51][62],
reservoir_weight[51][63],
reservoir_weight[51][64],
reservoir_weight[51][65],
reservoir_weight[51][66],
reservoir_weight[51][67],
reservoir_weight[51][68],
reservoir_weight[51][69],
reservoir_weight[51][70],
reservoir_weight[51][71],
reservoir_weight[51][72],
reservoir_weight[51][73],
reservoir_weight[51][74],
reservoir_weight[51][75],
reservoir_weight[51][76],
reservoir_weight[51][77],
reservoir_weight[51][78],
reservoir_weight[51][79],
reservoir_weight[51][80],
reservoir_weight[51][81],
reservoir_weight[51][82],
reservoir_weight[51][83],
reservoir_weight[51][84],
reservoir_weight[51][85],
reservoir_weight[51][86],
reservoir_weight[51][87],
reservoir_weight[51][88],
reservoir_weight[51][89],
reservoir_weight[51][90],
reservoir_weight[51][91],
reservoir_weight[51][92],
reservoir_weight[51][93],
reservoir_weight[51][94],
reservoir_weight[51][95],
reservoir_weight[51][96],
reservoir_weight[51][97],
reservoir_weight[51][98],
reservoir_weight[51][99],
reservoir_weight[51][100],
reservoir_weight[51][101],
reservoir_weight[51][102],
reservoir_weight[51][103],
reservoir_weight[51][104],
reservoir_weight[51][105],
reservoir_weight[51][106],
reservoir_weight[51][107],
reservoir_weight[51][108],
reservoir_weight[51][109],
reservoir_weight[51][110],
reservoir_weight[51][111],
reservoir_weight[51][112],
reservoir_weight[51][113],
reservoir_weight[51][114],
reservoir_weight[51][115],
reservoir_weight[51][116],
reservoir_weight[51][117],
reservoir_weight[51][118],
reservoir_weight[51][119],
reservoir_weight[51][120],
reservoir_weight[51][121],
reservoir_weight[51][122],
reservoir_weight[51][123],
reservoir_weight[51][124],
reservoir_weight[51][125],
reservoir_weight[51][126],
reservoir_weight[51][127],
reservoir_weight[51][128],
reservoir_weight[51][129],
reservoir_weight[51][130],
reservoir_weight[51][131],
reservoir_weight[51][132],
reservoir_weight[51][133],
reservoir_weight[51][134],
reservoir_weight[51][135],
reservoir_weight[51][136],
reservoir_weight[51][137],
reservoir_weight[51][138],
reservoir_weight[51][139],
reservoir_weight[51][140],
reservoir_weight[51][141],
reservoir_weight[51][142],
reservoir_weight[51][143],
reservoir_weight[51][144],
reservoir_weight[51][145],
reservoir_weight[51][146],
reservoir_weight[51][147],
reservoir_weight[51][148],
reservoir_weight[51][149],
reservoir_weight[51][150],
reservoir_weight[51][151],
reservoir_weight[51][152],
reservoir_weight[51][153],
reservoir_weight[51][154],
reservoir_weight[51][155],
reservoir_weight[51][156],
reservoir_weight[51][157],
reservoir_weight[51][158],
reservoir_weight[51][159],
reservoir_weight[51][160],
reservoir_weight[51][161],
reservoir_weight[51][162],
reservoir_weight[51][163],
reservoir_weight[51][164],
reservoir_weight[51][165],
reservoir_weight[51][166],
reservoir_weight[51][167],
reservoir_weight[51][168],
reservoir_weight[51][169],
reservoir_weight[51][170],
reservoir_weight[51][171],
reservoir_weight[51][172],
reservoir_weight[51][173],
reservoir_weight[51][174],
reservoir_weight[51][175],
reservoir_weight[51][176],
reservoir_weight[51][177],
reservoir_weight[51][178],
reservoir_weight[51][179],
reservoir_weight[51][180],
reservoir_weight[51][181],
reservoir_weight[51][182],
reservoir_weight[51][183],
reservoir_weight[51][184],
reservoir_weight[51][185],
reservoir_weight[51][186],
reservoir_weight[51][187],
reservoir_weight[51][188],
reservoir_weight[51][189],
reservoir_weight[51][190],
reservoir_weight[51][191],
reservoir_weight[51][192],
reservoir_weight[51][193],
reservoir_weight[51][194],
reservoir_weight[51][195],
reservoir_weight[51][196],
reservoir_weight[51][197],
reservoir_weight[51][198],
reservoir_weight[51][199]
},
{reservoir_weight[52][0],
reservoir_weight[52][1],
reservoir_weight[52][2],
reservoir_weight[52][3],
reservoir_weight[52][4],
reservoir_weight[52][5],
reservoir_weight[52][6],
reservoir_weight[52][7],
reservoir_weight[52][8],
reservoir_weight[52][9],
reservoir_weight[52][10],
reservoir_weight[52][11],
reservoir_weight[52][12],
reservoir_weight[52][13],
reservoir_weight[52][14],
reservoir_weight[52][15],
reservoir_weight[52][16],
reservoir_weight[52][17],
reservoir_weight[52][18],
reservoir_weight[52][19],
reservoir_weight[52][20],
reservoir_weight[52][21],
reservoir_weight[52][22],
reservoir_weight[52][23],
reservoir_weight[52][24],
reservoir_weight[52][25],
reservoir_weight[52][26],
reservoir_weight[52][27],
reservoir_weight[52][28],
reservoir_weight[52][29],
reservoir_weight[52][30],
reservoir_weight[52][31],
reservoir_weight[52][32],
reservoir_weight[52][33],
reservoir_weight[52][34],
reservoir_weight[52][35],
reservoir_weight[52][36],
reservoir_weight[52][37],
reservoir_weight[52][38],
reservoir_weight[52][39],
reservoir_weight[52][40],
reservoir_weight[52][41],
reservoir_weight[52][42],
reservoir_weight[52][43],
reservoir_weight[52][44],
reservoir_weight[52][45],
reservoir_weight[52][46],
reservoir_weight[52][47],
reservoir_weight[52][48],
reservoir_weight[52][49],
reservoir_weight[52][50],
reservoir_weight[52][51],
reservoir_weight[52][52],
reservoir_weight[52][53],
reservoir_weight[52][54],
reservoir_weight[52][55],
reservoir_weight[52][56],
reservoir_weight[52][57],
reservoir_weight[52][58],
reservoir_weight[52][59],
reservoir_weight[52][60],
reservoir_weight[52][61],
reservoir_weight[52][62],
reservoir_weight[52][63],
reservoir_weight[52][64],
reservoir_weight[52][65],
reservoir_weight[52][66],
reservoir_weight[52][67],
reservoir_weight[52][68],
reservoir_weight[52][69],
reservoir_weight[52][70],
reservoir_weight[52][71],
reservoir_weight[52][72],
reservoir_weight[52][73],
reservoir_weight[52][74],
reservoir_weight[52][75],
reservoir_weight[52][76],
reservoir_weight[52][77],
reservoir_weight[52][78],
reservoir_weight[52][79],
reservoir_weight[52][80],
reservoir_weight[52][81],
reservoir_weight[52][82],
reservoir_weight[52][83],
reservoir_weight[52][84],
reservoir_weight[52][85],
reservoir_weight[52][86],
reservoir_weight[52][87],
reservoir_weight[52][88],
reservoir_weight[52][89],
reservoir_weight[52][90],
reservoir_weight[52][91],
reservoir_weight[52][92],
reservoir_weight[52][93],
reservoir_weight[52][94],
reservoir_weight[52][95],
reservoir_weight[52][96],
reservoir_weight[52][97],
reservoir_weight[52][98],
reservoir_weight[52][99],
reservoir_weight[52][100],
reservoir_weight[52][101],
reservoir_weight[52][102],
reservoir_weight[52][103],
reservoir_weight[52][104],
reservoir_weight[52][105],
reservoir_weight[52][106],
reservoir_weight[52][107],
reservoir_weight[52][108],
reservoir_weight[52][109],
reservoir_weight[52][110],
reservoir_weight[52][111],
reservoir_weight[52][112],
reservoir_weight[52][113],
reservoir_weight[52][114],
reservoir_weight[52][115],
reservoir_weight[52][116],
reservoir_weight[52][117],
reservoir_weight[52][118],
reservoir_weight[52][119],
reservoir_weight[52][120],
reservoir_weight[52][121],
reservoir_weight[52][122],
reservoir_weight[52][123],
reservoir_weight[52][124],
reservoir_weight[52][125],
reservoir_weight[52][126],
reservoir_weight[52][127],
reservoir_weight[52][128],
reservoir_weight[52][129],
reservoir_weight[52][130],
reservoir_weight[52][131],
reservoir_weight[52][132],
reservoir_weight[52][133],
reservoir_weight[52][134],
reservoir_weight[52][135],
reservoir_weight[52][136],
reservoir_weight[52][137],
reservoir_weight[52][138],
reservoir_weight[52][139],
reservoir_weight[52][140],
reservoir_weight[52][141],
reservoir_weight[52][142],
reservoir_weight[52][143],
reservoir_weight[52][144],
reservoir_weight[52][145],
reservoir_weight[52][146],
reservoir_weight[52][147],
reservoir_weight[52][148],
reservoir_weight[52][149],
reservoir_weight[52][150],
reservoir_weight[52][151],
reservoir_weight[52][152],
reservoir_weight[52][153],
reservoir_weight[52][154],
reservoir_weight[52][155],
reservoir_weight[52][156],
reservoir_weight[52][157],
reservoir_weight[52][158],
reservoir_weight[52][159],
reservoir_weight[52][160],
reservoir_weight[52][161],
reservoir_weight[52][162],
reservoir_weight[52][163],
reservoir_weight[52][164],
reservoir_weight[52][165],
reservoir_weight[52][166],
reservoir_weight[52][167],
reservoir_weight[52][168],
reservoir_weight[52][169],
reservoir_weight[52][170],
reservoir_weight[52][171],
reservoir_weight[52][172],
reservoir_weight[52][173],
reservoir_weight[52][174],
reservoir_weight[52][175],
reservoir_weight[52][176],
reservoir_weight[52][177],
reservoir_weight[52][178],
reservoir_weight[52][179],
reservoir_weight[52][180],
reservoir_weight[52][181],
reservoir_weight[52][182],
reservoir_weight[52][183],
reservoir_weight[52][184],
reservoir_weight[52][185],
reservoir_weight[52][186],
reservoir_weight[52][187],
reservoir_weight[52][188],
reservoir_weight[52][189],
reservoir_weight[52][190],
reservoir_weight[52][191],
reservoir_weight[52][192],
reservoir_weight[52][193],
reservoir_weight[52][194],
reservoir_weight[52][195],
reservoir_weight[52][196],
reservoir_weight[52][197],
reservoir_weight[52][198],
reservoir_weight[52][199]
},
{reservoir_weight[53][0],
reservoir_weight[53][1],
reservoir_weight[53][2],
reservoir_weight[53][3],
reservoir_weight[53][4],
reservoir_weight[53][5],
reservoir_weight[53][6],
reservoir_weight[53][7],
reservoir_weight[53][8],
reservoir_weight[53][9],
reservoir_weight[53][10],
reservoir_weight[53][11],
reservoir_weight[53][12],
reservoir_weight[53][13],
reservoir_weight[53][14],
reservoir_weight[53][15],
reservoir_weight[53][16],
reservoir_weight[53][17],
reservoir_weight[53][18],
reservoir_weight[53][19],
reservoir_weight[53][20],
reservoir_weight[53][21],
reservoir_weight[53][22],
reservoir_weight[53][23],
reservoir_weight[53][24],
reservoir_weight[53][25],
reservoir_weight[53][26],
reservoir_weight[53][27],
reservoir_weight[53][28],
reservoir_weight[53][29],
reservoir_weight[53][30],
reservoir_weight[53][31],
reservoir_weight[53][32],
reservoir_weight[53][33],
reservoir_weight[53][34],
reservoir_weight[53][35],
reservoir_weight[53][36],
reservoir_weight[53][37],
reservoir_weight[53][38],
reservoir_weight[53][39],
reservoir_weight[53][40],
reservoir_weight[53][41],
reservoir_weight[53][42],
reservoir_weight[53][43],
reservoir_weight[53][44],
reservoir_weight[53][45],
reservoir_weight[53][46],
reservoir_weight[53][47],
reservoir_weight[53][48],
reservoir_weight[53][49],
reservoir_weight[53][50],
reservoir_weight[53][51],
reservoir_weight[53][52],
reservoir_weight[53][53],
reservoir_weight[53][54],
reservoir_weight[53][55],
reservoir_weight[53][56],
reservoir_weight[53][57],
reservoir_weight[53][58],
reservoir_weight[53][59],
reservoir_weight[53][60],
reservoir_weight[53][61],
reservoir_weight[53][62],
reservoir_weight[53][63],
reservoir_weight[53][64],
reservoir_weight[53][65],
reservoir_weight[53][66],
reservoir_weight[53][67],
reservoir_weight[53][68],
reservoir_weight[53][69],
reservoir_weight[53][70],
reservoir_weight[53][71],
reservoir_weight[53][72],
reservoir_weight[53][73],
reservoir_weight[53][74],
reservoir_weight[53][75],
reservoir_weight[53][76],
reservoir_weight[53][77],
reservoir_weight[53][78],
reservoir_weight[53][79],
reservoir_weight[53][80],
reservoir_weight[53][81],
reservoir_weight[53][82],
reservoir_weight[53][83],
reservoir_weight[53][84],
reservoir_weight[53][85],
reservoir_weight[53][86],
reservoir_weight[53][87],
reservoir_weight[53][88],
reservoir_weight[53][89],
reservoir_weight[53][90],
reservoir_weight[53][91],
reservoir_weight[53][92],
reservoir_weight[53][93],
reservoir_weight[53][94],
reservoir_weight[53][95],
reservoir_weight[53][96],
reservoir_weight[53][97],
reservoir_weight[53][98],
reservoir_weight[53][99],
reservoir_weight[53][100],
reservoir_weight[53][101],
reservoir_weight[53][102],
reservoir_weight[53][103],
reservoir_weight[53][104],
reservoir_weight[53][105],
reservoir_weight[53][106],
reservoir_weight[53][107],
reservoir_weight[53][108],
reservoir_weight[53][109],
reservoir_weight[53][110],
reservoir_weight[53][111],
reservoir_weight[53][112],
reservoir_weight[53][113],
reservoir_weight[53][114],
reservoir_weight[53][115],
reservoir_weight[53][116],
reservoir_weight[53][117],
reservoir_weight[53][118],
reservoir_weight[53][119],
reservoir_weight[53][120],
reservoir_weight[53][121],
reservoir_weight[53][122],
reservoir_weight[53][123],
reservoir_weight[53][124],
reservoir_weight[53][125],
reservoir_weight[53][126],
reservoir_weight[53][127],
reservoir_weight[53][128],
reservoir_weight[53][129],
reservoir_weight[53][130],
reservoir_weight[53][131],
reservoir_weight[53][132],
reservoir_weight[53][133],
reservoir_weight[53][134],
reservoir_weight[53][135],
reservoir_weight[53][136],
reservoir_weight[53][137],
reservoir_weight[53][138],
reservoir_weight[53][139],
reservoir_weight[53][140],
reservoir_weight[53][141],
reservoir_weight[53][142],
reservoir_weight[53][143],
reservoir_weight[53][144],
reservoir_weight[53][145],
reservoir_weight[53][146],
reservoir_weight[53][147],
reservoir_weight[53][148],
reservoir_weight[53][149],
reservoir_weight[53][150],
reservoir_weight[53][151],
reservoir_weight[53][152],
reservoir_weight[53][153],
reservoir_weight[53][154],
reservoir_weight[53][155],
reservoir_weight[53][156],
reservoir_weight[53][157],
reservoir_weight[53][158],
reservoir_weight[53][159],
reservoir_weight[53][160],
reservoir_weight[53][161],
reservoir_weight[53][162],
reservoir_weight[53][163],
reservoir_weight[53][164],
reservoir_weight[53][165],
reservoir_weight[53][166],
reservoir_weight[53][167],
reservoir_weight[53][168],
reservoir_weight[53][169],
reservoir_weight[53][170],
reservoir_weight[53][171],
reservoir_weight[53][172],
reservoir_weight[53][173],
reservoir_weight[53][174],
reservoir_weight[53][175],
reservoir_weight[53][176],
reservoir_weight[53][177],
reservoir_weight[53][178],
reservoir_weight[53][179],
reservoir_weight[53][180],
reservoir_weight[53][181],
reservoir_weight[53][182],
reservoir_weight[53][183],
reservoir_weight[53][184],
reservoir_weight[53][185],
reservoir_weight[53][186],
reservoir_weight[53][187],
reservoir_weight[53][188],
reservoir_weight[53][189],
reservoir_weight[53][190],
reservoir_weight[53][191],
reservoir_weight[53][192],
reservoir_weight[53][193],
reservoir_weight[53][194],
reservoir_weight[53][195],
reservoir_weight[53][196],
reservoir_weight[53][197],
reservoir_weight[53][198],
reservoir_weight[53][199]
},
{reservoir_weight[54][0],
reservoir_weight[54][1],
reservoir_weight[54][2],
reservoir_weight[54][3],
reservoir_weight[54][4],
reservoir_weight[54][5],
reservoir_weight[54][6],
reservoir_weight[54][7],
reservoir_weight[54][8],
reservoir_weight[54][9],
reservoir_weight[54][10],
reservoir_weight[54][11],
reservoir_weight[54][12],
reservoir_weight[54][13],
reservoir_weight[54][14],
reservoir_weight[54][15],
reservoir_weight[54][16],
reservoir_weight[54][17],
reservoir_weight[54][18],
reservoir_weight[54][19],
reservoir_weight[54][20],
reservoir_weight[54][21],
reservoir_weight[54][22],
reservoir_weight[54][23],
reservoir_weight[54][24],
reservoir_weight[54][25],
reservoir_weight[54][26],
reservoir_weight[54][27],
reservoir_weight[54][28],
reservoir_weight[54][29],
reservoir_weight[54][30],
reservoir_weight[54][31],
reservoir_weight[54][32],
reservoir_weight[54][33],
reservoir_weight[54][34],
reservoir_weight[54][35],
reservoir_weight[54][36],
reservoir_weight[54][37],
reservoir_weight[54][38],
reservoir_weight[54][39],
reservoir_weight[54][40],
reservoir_weight[54][41],
reservoir_weight[54][42],
reservoir_weight[54][43],
reservoir_weight[54][44],
reservoir_weight[54][45],
reservoir_weight[54][46],
reservoir_weight[54][47],
reservoir_weight[54][48],
reservoir_weight[54][49],
reservoir_weight[54][50],
reservoir_weight[54][51],
reservoir_weight[54][52],
reservoir_weight[54][53],
reservoir_weight[54][54],
reservoir_weight[54][55],
reservoir_weight[54][56],
reservoir_weight[54][57],
reservoir_weight[54][58],
reservoir_weight[54][59],
reservoir_weight[54][60],
reservoir_weight[54][61],
reservoir_weight[54][62],
reservoir_weight[54][63],
reservoir_weight[54][64],
reservoir_weight[54][65],
reservoir_weight[54][66],
reservoir_weight[54][67],
reservoir_weight[54][68],
reservoir_weight[54][69],
reservoir_weight[54][70],
reservoir_weight[54][71],
reservoir_weight[54][72],
reservoir_weight[54][73],
reservoir_weight[54][74],
reservoir_weight[54][75],
reservoir_weight[54][76],
reservoir_weight[54][77],
reservoir_weight[54][78],
reservoir_weight[54][79],
reservoir_weight[54][80],
reservoir_weight[54][81],
reservoir_weight[54][82],
reservoir_weight[54][83],
reservoir_weight[54][84],
reservoir_weight[54][85],
reservoir_weight[54][86],
reservoir_weight[54][87],
reservoir_weight[54][88],
reservoir_weight[54][89],
reservoir_weight[54][90],
reservoir_weight[54][91],
reservoir_weight[54][92],
reservoir_weight[54][93],
reservoir_weight[54][94],
reservoir_weight[54][95],
reservoir_weight[54][96],
reservoir_weight[54][97],
reservoir_weight[54][98],
reservoir_weight[54][99],
reservoir_weight[54][100],
reservoir_weight[54][101],
reservoir_weight[54][102],
reservoir_weight[54][103],
reservoir_weight[54][104],
reservoir_weight[54][105],
reservoir_weight[54][106],
reservoir_weight[54][107],
reservoir_weight[54][108],
reservoir_weight[54][109],
reservoir_weight[54][110],
reservoir_weight[54][111],
reservoir_weight[54][112],
reservoir_weight[54][113],
reservoir_weight[54][114],
reservoir_weight[54][115],
reservoir_weight[54][116],
reservoir_weight[54][117],
reservoir_weight[54][118],
reservoir_weight[54][119],
reservoir_weight[54][120],
reservoir_weight[54][121],
reservoir_weight[54][122],
reservoir_weight[54][123],
reservoir_weight[54][124],
reservoir_weight[54][125],
reservoir_weight[54][126],
reservoir_weight[54][127],
reservoir_weight[54][128],
reservoir_weight[54][129],
reservoir_weight[54][130],
reservoir_weight[54][131],
reservoir_weight[54][132],
reservoir_weight[54][133],
reservoir_weight[54][134],
reservoir_weight[54][135],
reservoir_weight[54][136],
reservoir_weight[54][137],
reservoir_weight[54][138],
reservoir_weight[54][139],
reservoir_weight[54][140],
reservoir_weight[54][141],
reservoir_weight[54][142],
reservoir_weight[54][143],
reservoir_weight[54][144],
reservoir_weight[54][145],
reservoir_weight[54][146],
reservoir_weight[54][147],
reservoir_weight[54][148],
reservoir_weight[54][149],
reservoir_weight[54][150],
reservoir_weight[54][151],
reservoir_weight[54][152],
reservoir_weight[54][153],
reservoir_weight[54][154],
reservoir_weight[54][155],
reservoir_weight[54][156],
reservoir_weight[54][157],
reservoir_weight[54][158],
reservoir_weight[54][159],
reservoir_weight[54][160],
reservoir_weight[54][161],
reservoir_weight[54][162],
reservoir_weight[54][163],
reservoir_weight[54][164],
reservoir_weight[54][165],
reservoir_weight[54][166],
reservoir_weight[54][167],
reservoir_weight[54][168],
reservoir_weight[54][169],
reservoir_weight[54][170],
reservoir_weight[54][171],
reservoir_weight[54][172],
reservoir_weight[54][173],
reservoir_weight[54][174],
reservoir_weight[54][175],
reservoir_weight[54][176],
reservoir_weight[54][177],
reservoir_weight[54][178],
reservoir_weight[54][179],
reservoir_weight[54][180],
reservoir_weight[54][181],
reservoir_weight[54][182],
reservoir_weight[54][183],
reservoir_weight[54][184],
reservoir_weight[54][185],
reservoir_weight[54][186],
reservoir_weight[54][187],
reservoir_weight[54][188],
reservoir_weight[54][189],
reservoir_weight[54][190],
reservoir_weight[54][191],
reservoir_weight[54][192],
reservoir_weight[54][193],
reservoir_weight[54][194],
reservoir_weight[54][195],
reservoir_weight[54][196],
reservoir_weight[54][197],
reservoir_weight[54][198],
reservoir_weight[54][199]
},
{reservoir_weight[55][0],
reservoir_weight[55][1],
reservoir_weight[55][2],
reservoir_weight[55][3],
reservoir_weight[55][4],
reservoir_weight[55][5],
reservoir_weight[55][6],
reservoir_weight[55][7],
reservoir_weight[55][8],
reservoir_weight[55][9],
reservoir_weight[55][10],
reservoir_weight[55][11],
reservoir_weight[55][12],
reservoir_weight[55][13],
reservoir_weight[55][14],
reservoir_weight[55][15],
reservoir_weight[55][16],
reservoir_weight[55][17],
reservoir_weight[55][18],
reservoir_weight[55][19],
reservoir_weight[55][20],
reservoir_weight[55][21],
reservoir_weight[55][22],
reservoir_weight[55][23],
reservoir_weight[55][24],
reservoir_weight[55][25],
reservoir_weight[55][26],
reservoir_weight[55][27],
reservoir_weight[55][28],
reservoir_weight[55][29],
reservoir_weight[55][30],
reservoir_weight[55][31],
reservoir_weight[55][32],
reservoir_weight[55][33],
reservoir_weight[55][34],
reservoir_weight[55][35],
reservoir_weight[55][36],
reservoir_weight[55][37],
reservoir_weight[55][38],
reservoir_weight[55][39],
reservoir_weight[55][40],
reservoir_weight[55][41],
reservoir_weight[55][42],
reservoir_weight[55][43],
reservoir_weight[55][44],
reservoir_weight[55][45],
reservoir_weight[55][46],
reservoir_weight[55][47],
reservoir_weight[55][48],
reservoir_weight[55][49],
reservoir_weight[55][50],
reservoir_weight[55][51],
reservoir_weight[55][52],
reservoir_weight[55][53],
reservoir_weight[55][54],
reservoir_weight[55][55],
reservoir_weight[55][56],
reservoir_weight[55][57],
reservoir_weight[55][58],
reservoir_weight[55][59],
reservoir_weight[55][60],
reservoir_weight[55][61],
reservoir_weight[55][62],
reservoir_weight[55][63],
reservoir_weight[55][64],
reservoir_weight[55][65],
reservoir_weight[55][66],
reservoir_weight[55][67],
reservoir_weight[55][68],
reservoir_weight[55][69],
reservoir_weight[55][70],
reservoir_weight[55][71],
reservoir_weight[55][72],
reservoir_weight[55][73],
reservoir_weight[55][74],
reservoir_weight[55][75],
reservoir_weight[55][76],
reservoir_weight[55][77],
reservoir_weight[55][78],
reservoir_weight[55][79],
reservoir_weight[55][80],
reservoir_weight[55][81],
reservoir_weight[55][82],
reservoir_weight[55][83],
reservoir_weight[55][84],
reservoir_weight[55][85],
reservoir_weight[55][86],
reservoir_weight[55][87],
reservoir_weight[55][88],
reservoir_weight[55][89],
reservoir_weight[55][90],
reservoir_weight[55][91],
reservoir_weight[55][92],
reservoir_weight[55][93],
reservoir_weight[55][94],
reservoir_weight[55][95],
reservoir_weight[55][96],
reservoir_weight[55][97],
reservoir_weight[55][98],
reservoir_weight[55][99],
reservoir_weight[55][100],
reservoir_weight[55][101],
reservoir_weight[55][102],
reservoir_weight[55][103],
reservoir_weight[55][104],
reservoir_weight[55][105],
reservoir_weight[55][106],
reservoir_weight[55][107],
reservoir_weight[55][108],
reservoir_weight[55][109],
reservoir_weight[55][110],
reservoir_weight[55][111],
reservoir_weight[55][112],
reservoir_weight[55][113],
reservoir_weight[55][114],
reservoir_weight[55][115],
reservoir_weight[55][116],
reservoir_weight[55][117],
reservoir_weight[55][118],
reservoir_weight[55][119],
reservoir_weight[55][120],
reservoir_weight[55][121],
reservoir_weight[55][122],
reservoir_weight[55][123],
reservoir_weight[55][124],
reservoir_weight[55][125],
reservoir_weight[55][126],
reservoir_weight[55][127],
reservoir_weight[55][128],
reservoir_weight[55][129],
reservoir_weight[55][130],
reservoir_weight[55][131],
reservoir_weight[55][132],
reservoir_weight[55][133],
reservoir_weight[55][134],
reservoir_weight[55][135],
reservoir_weight[55][136],
reservoir_weight[55][137],
reservoir_weight[55][138],
reservoir_weight[55][139],
reservoir_weight[55][140],
reservoir_weight[55][141],
reservoir_weight[55][142],
reservoir_weight[55][143],
reservoir_weight[55][144],
reservoir_weight[55][145],
reservoir_weight[55][146],
reservoir_weight[55][147],
reservoir_weight[55][148],
reservoir_weight[55][149],
reservoir_weight[55][150],
reservoir_weight[55][151],
reservoir_weight[55][152],
reservoir_weight[55][153],
reservoir_weight[55][154],
reservoir_weight[55][155],
reservoir_weight[55][156],
reservoir_weight[55][157],
reservoir_weight[55][158],
reservoir_weight[55][159],
reservoir_weight[55][160],
reservoir_weight[55][161],
reservoir_weight[55][162],
reservoir_weight[55][163],
reservoir_weight[55][164],
reservoir_weight[55][165],
reservoir_weight[55][166],
reservoir_weight[55][167],
reservoir_weight[55][168],
reservoir_weight[55][169],
reservoir_weight[55][170],
reservoir_weight[55][171],
reservoir_weight[55][172],
reservoir_weight[55][173],
reservoir_weight[55][174],
reservoir_weight[55][175],
reservoir_weight[55][176],
reservoir_weight[55][177],
reservoir_weight[55][178],
reservoir_weight[55][179],
reservoir_weight[55][180],
reservoir_weight[55][181],
reservoir_weight[55][182],
reservoir_weight[55][183],
reservoir_weight[55][184],
reservoir_weight[55][185],
reservoir_weight[55][186],
reservoir_weight[55][187],
reservoir_weight[55][188],
reservoir_weight[55][189],
reservoir_weight[55][190],
reservoir_weight[55][191],
reservoir_weight[55][192],
reservoir_weight[55][193],
reservoir_weight[55][194],
reservoir_weight[55][195],
reservoir_weight[55][196],
reservoir_weight[55][197],
reservoir_weight[55][198],
reservoir_weight[55][199]
},
{reservoir_weight[56][0],
reservoir_weight[56][1],
reservoir_weight[56][2],
reservoir_weight[56][3],
reservoir_weight[56][4],
reservoir_weight[56][5],
reservoir_weight[56][6],
reservoir_weight[56][7],
reservoir_weight[56][8],
reservoir_weight[56][9],
reservoir_weight[56][10],
reservoir_weight[56][11],
reservoir_weight[56][12],
reservoir_weight[56][13],
reservoir_weight[56][14],
reservoir_weight[56][15],
reservoir_weight[56][16],
reservoir_weight[56][17],
reservoir_weight[56][18],
reservoir_weight[56][19],
reservoir_weight[56][20],
reservoir_weight[56][21],
reservoir_weight[56][22],
reservoir_weight[56][23],
reservoir_weight[56][24],
reservoir_weight[56][25],
reservoir_weight[56][26],
reservoir_weight[56][27],
reservoir_weight[56][28],
reservoir_weight[56][29],
reservoir_weight[56][30],
reservoir_weight[56][31],
reservoir_weight[56][32],
reservoir_weight[56][33],
reservoir_weight[56][34],
reservoir_weight[56][35],
reservoir_weight[56][36],
reservoir_weight[56][37],
reservoir_weight[56][38],
reservoir_weight[56][39],
reservoir_weight[56][40],
reservoir_weight[56][41],
reservoir_weight[56][42],
reservoir_weight[56][43],
reservoir_weight[56][44],
reservoir_weight[56][45],
reservoir_weight[56][46],
reservoir_weight[56][47],
reservoir_weight[56][48],
reservoir_weight[56][49],
reservoir_weight[56][50],
reservoir_weight[56][51],
reservoir_weight[56][52],
reservoir_weight[56][53],
reservoir_weight[56][54],
reservoir_weight[56][55],
reservoir_weight[56][56],
reservoir_weight[56][57],
reservoir_weight[56][58],
reservoir_weight[56][59],
reservoir_weight[56][60],
reservoir_weight[56][61],
reservoir_weight[56][62],
reservoir_weight[56][63],
reservoir_weight[56][64],
reservoir_weight[56][65],
reservoir_weight[56][66],
reservoir_weight[56][67],
reservoir_weight[56][68],
reservoir_weight[56][69],
reservoir_weight[56][70],
reservoir_weight[56][71],
reservoir_weight[56][72],
reservoir_weight[56][73],
reservoir_weight[56][74],
reservoir_weight[56][75],
reservoir_weight[56][76],
reservoir_weight[56][77],
reservoir_weight[56][78],
reservoir_weight[56][79],
reservoir_weight[56][80],
reservoir_weight[56][81],
reservoir_weight[56][82],
reservoir_weight[56][83],
reservoir_weight[56][84],
reservoir_weight[56][85],
reservoir_weight[56][86],
reservoir_weight[56][87],
reservoir_weight[56][88],
reservoir_weight[56][89],
reservoir_weight[56][90],
reservoir_weight[56][91],
reservoir_weight[56][92],
reservoir_weight[56][93],
reservoir_weight[56][94],
reservoir_weight[56][95],
reservoir_weight[56][96],
reservoir_weight[56][97],
reservoir_weight[56][98],
reservoir_weight[56][99],
reservoir_weight[56][100],
reservoir_weight[56][101],
reservoir_weight[56][102],
reservoir_weight[56][103],
reservoir_weight[56][104],
reservoir_weight[56][105],
reservoir_weight[56][106],
reservoir_weight[56][107],
reservoir_weight[56][108],
reservoir_weight[56][109],
reservoir_weight[56][110],
reservoir_weight[56][111],
reservoir_weight[56][112],
reservoir_weight[56][113],
reservoir_weight[56][114],
reservoir_weight[56][115],
reservoir_weight[56][116],
reservoir_weight[56][117],
reservoir_weight[56][118],
reservoir_weight[56][119],
reservoir_weight[56][120],
reservoir_weight[56][121],
reservoir_weight[56][122],
reservoir_weight[56][123],
reservoir_weight[56][124],
reservoir_weight[56][125],
reservoir_weight[56][126],
reservoir_weight[56][127],
reservoir_weight[56][128],
reservoir_weight[56][129],
reservoir_weight[56][130],
reservoir_weight[56][131],
reservoir_weight[56][132],
reservoir_weight[56][133],
reservoir_weight[56][134],
reservoir_weight[56][135],
reservoir_weight[56][136],
reservoir_weight[56][137],
reservoir_weight[56][138],
reservoir_weight[56][139],
reservoir_weight[56][140],
reservoir_weight[56][141],
reservoir_weight[56][142],
reservoir_weight[56][143],
reservoir_weight[56][144],
reservoir_weight[56][145],
reservoir_weight[56][146],
reservoir_weight[56][147],
reservoir_weight[56][148],
reservoir_weight[56][149],
reservoir_weight[56][150],
reservoir_weight[56][151],
reservoir_weight[56][152],
reservoir_weight[56][153],
reservoir_weight[56][154],
reservoir_weight[56][155],
reservoir_weight[56][156],
reservoir_weight[56][157],
reservoir_weight[56][158],
reservoir_weight[56][159],
reservoir_weight[56][160],
reservoir_weight[56][161],
reservoir_weight[56][162],
reservoir_weight[56][163],
reservoir_weight[56][164],
reservoir_weight[56][165],
reservoir_weight[56][166],
reservoir_weight[56][167],
reservoir_weight[56][168],
reservoir_weight[56][169],
reservoir_weight[56][170],
reservoir_weight[56][171],
reservoir_weight[56][172],
reservoir_weight[56][173],
reservoir_weight[56][174],
reservoir_weight[56][175],
reservoir_weight[56][176],
reservoir_weight[56][177],
reservoir_weight[56][178],
reservoir_weight[56][179],
reservoir_weight[56][180],
reservoir_weight[56][181],
reservoir_weight[56][182],
reservoir_weight[56][183],
reservoir_weight[56][184],
reservoir_weight[56][185],
reservoir_weight[56][186],
reservoir_weight[56][187],
reservoir_weight[56][188],
reservoir_weight[56][189],
reservoir_weight[56][190],
reservoir_weight[56][191],
reservoir_weight[56][192],
reservoir_weight[56][193],
reservoir_weight[56][194],
reservoir_weight[56][195],
reservoir_weight[56][196],
reservoir_weight[56][197],
reservoir_weight[56][198],
reservoir_weight[56][199]
},
{reservoir_weight[57][0],
reservoir_weight[57][1],
reservoir_weight[57][2],
reservoir_weight[57][3],
reservoir_weight[57][4],
reservoir_weight[57][5],
reservoir_weight[57][6],
reservoir_weight[57][7],
reservoir_weight[57][8],
reservoir_weight[57][9],
reservoir_weight[57][10],
reservoir_weight[57][11],
reservoir_weight[57][12],
reservoir_weight[57][13],
reservoir_weight[57][14],
reservoir_weight[57][15],
reservoir_weight[57][16],
reservoir_weight[57][17],
reservoir_weight[57][18],
reservoir_weight[57][19],
reservoir_weight[57][20],
reservoir_weight[57][21],
reservoir_weight[57][22],
reservoir_weight[57][23],
reservoir_weight[57][24],
reservoir_weight[57][25],
reservoir_weight[57][26],
reservoir_weight[57][27],
reservoir_weight[57][28],
reservoir_weight[57][29],
reservoir_weight[57][30],
reservoir_weight[57][31],
reservoir_weight[57][32],
reservoir_weight[57][33],
reservoir_weight[57][34],
reservoir_weight[57][35],
reservoir_weight[57][36],
reservoir_weight[57][37],
reservoir_weight[57][38],
reservoir_weight[57][39],
reservoir_weight[57][40],
reservoir_weight[57][41],
reservoir_weight[57][42],
reservoir_weight[57][43],
reservoir_weight[57][44],
reservoir_weight[57][45],
reservoir_weight[57][46],
reservoir_weight[57][47],
reservoir_weight[57][48],
reservoir_weight[57][49],
reservoir_weight[57][50],
reservoir_weight[57][51],
reservoir_weight[57][52],
reservoir_weight[57][53],
reservoir_weight[57][54],
reservoir_weight[57][55],
reservoir_weight[57][56],
reservoir_weight[57][57],
reservoir_weight[57][58],
reservoir_weight[57][59],
reservoir_weight[57][60],
reservoir_weight[57][61],
reservoir_weight[57][62],
reservoir_weight[57][63],
reservoir_weight[57][64],
reservoir_weight[57][65],
reservoir_weight[57][66],
reservoir_weight[57][67],
reservoir_weight[57][68],
reservoir_weight[57][69],
reservoir_weight[57][70],
reservoir_weight[57][71],
reservoir_weight[57][72],
reservoir_weight[57][73],
reservoir_weight[57][74],
reservoir_weight[57][75],
reservoir_weight[57][76],
reservoir_weight[57][77],
reservoir_weight[57][78],
reservoir_weight[57][79],
reservoir_weight[57][80],
reservoir_weight[57][81],
reservoir_weight[57][82],
reservoir_weight[57][83],
reservoir_weight[57][84],
reservoir_weight[57][85],
reservoir_weight[57][86],
reservoir_weight[57][87],
reservoir_weight[57][88],
reservoir_weight[57][89],
reservoir_weight[57][90],
reservoir_weight[57][91],
reservoir_weight[57][92],
reservoir_weight[57][93],
reservoir_weight[57][94],
reservoir_weight[57][95],
reservoir_weight[57][96],
reservoir_weight[57][97],
reservoir_weight[57][98],
reservoir_weight[57][99],
reservoir_weight[57][100],
reservoir_weight[57][101],
reservoir_weight[57][102],
reservoir_weight[57][103],
reservoir_weight[57][104],
reservoir_weight[57][105],
reservoir_weight[57][106],
reservoir_weight[57][107],
reservoir_weight[57][108],
reservoir_weight[57][109],
reservoir_weight[57][110],
reservoir_weight[57][111],
reservoir_weight[57][112],
reservoir_weight[57][113],
reservoir_weight[57][114],
reservoir_weight[57][115],
reservoir_weight[57][116],
reservoir_weight[57][117],
reservoir_weight[57][118],
reservoir_weight[57][119],
reservoir_weight[57][120],
reservoir_weight[57][121],
reservoir_weight[57][122],
reservoir_weight[57][123],
reservoir_weight[57][124],
reservoir_weight[57][125],
reservoir_weight[57][126],
reservoir_weight[57][127],
reservoir_weight[57][128],
reservoir_weight[57][129],
reservoir_weight[57][130],
reservoir_weight[57][131],
reservoir_weight[57][132],
reservoir_weight[57][133],
reservoir_weight[57][134],
reservoir_weight[57][135],
reservoir_weight[57][136],
reservoir_weight[57][137],
reservoir_weight[57][138],
reservoir_weight[57][139],
reservoir_weight[57][140],
reservoir_weight[57][141],
reservoir_weight[57][142],
reservoir_weight[57][143],
reservoir_weight[57][144],
reservoir_weight[57][145],
reservoir_weight[57][146],
reservoir_weight[57][147],
reservoir_weight[57][148],
reservoir_weight[57][149],
reservoir_weight[57][150],
reservoir_weight[57][151],
reservoir_weight[57][152],
reservoir_weight[57][153],
reservoir_weight[57][154],
reservoir_weight[57][155],
reservoir_weight[57][156],
reservoir_weight[57][157],
reservoir_weight[57][158],
reservoir_weight[57][159],
reservoir_weight[57][160],
reservoir_weight[57][161],
reservoir_weight[57][162],
reservoir_weight[57][163],
reservoir_weight[57][164],
reservoir_weight[57][165],
reservoir_weight[57][166],
reservoir_weight[57][167],
reservoir_weight[57][168],
reservoir_weight[57][169],
reservoir_weight[57][170],
reservoir_weight[57][171],
reservoir_weight[57][172],
reservoir_weight[57][173],
reservoir_weight[57][174],
reservoir_weight[57][175],
reservoir_weight[57][176],
reservoir_weight[57][177],
reservoir_weight[57][178],
reservoir_weight[57][179],
reservoir_weight[57][180],
reservoir_weight[57][181],
reservoir_weight[57][182],
reservoir_weight[57][183],
reservoir_weight[57][184],
reservoir_weight[57][185],
reservoir_weight[57][186],
reservoir_weight[57][187],
reservoir_weight[57][188],
reservoir_weight[57][189],
reservoir_weight[57][190],
reservoir_weight[57][191],
reservoir_weight[57][192],
reservoir_weight[57][193],
reservoir_weight[57][194],
reservoir_weight[57][195],
reservoir_weight[57][196],
reservoir_weight[57][197],
reservoir_weight[57][198],
reservoir_weight[57][199]
},
{reservoir_weight[58][0],
reservoir_weight[58][1],
reservoir_weight[58][2],
reservoir_weight[58][3],
reservoir_weight[58][4],
reservoir_weight[58][5],
reservoir_weight[58][6],
reservoir_weight[58][7],
reservoir_weight[58][8],
reservoir_weight[58][9],
reservoir_weight[58][10],
reservoir_weight[58][11],
reservoir_weight[58][12],
reservoir_weight[58][13],
reservoir_weight[58][14],
reservoir_weight[58][15],
reservoir_weight[58][16],
reservoir_weight[58][17],
reservoir_weight[58][18],
reservoir_weight[58][19],
reservoir_weight[58][20],
reservoir_weight[58][21],
reservoir_weight[58][22],
reservoir_weight[58][23],
reservoir_weight[58][24],
reservoir_weight[58][25],
reservoir_weight[58][26],
reservoir_weight[58][27],
reservoir_weight[58][28],
reservoir_weight[58][29],
reservoir_weight[58][30],
reservoir_weight[58][31],
reservoir_weight[58][32],
reservoir_weight[58][33],
reservoir_weight[58][34],
reservoir_weight[58][35],
reservoir_weight[58][36],
reservoir_weight[58][37],
reservoir_weight[58][38],
reservoir_weight[58][39],
reservoir_weight[58][40],
reservoir_weight[58][41],
reservoir_weight[58][42],
reservoir_weight[58][43],
reservoir_weight[58][44],
reservoir_weight[58][45],
reservoir_weight[58][46],
reservoir_weight[58][47],
reservoir_weight[58][48],
reservoir_weight[58][49],
reservoir_weight[58][50],
reservoir_weight[58][51],
reservoir_weight[58][52],
reservoir_weight[58][53],
reservoir_weight[58][54],
reservoir_weight[58][55],
reservoir_weight[58][56],
reservoir_weight[58][57],
reservoir_weight[58][58],
reservoir_weight[58][59],
reservoir_weight[58][60],
reservoir_weight[58][61],
reservoir_weight[58][62],
reservoir_weight[58][63],
reservoir_weight[58][64],
reservoir_weight[58][65],
reservoir_weight[58][66],
reservoir_weight[58][67],
reservoir_weight[58][68],
reservoir_weight[58][69],
reservoir_weight[58][70],
reservoir_weight[58][71],
reservoir_weight[58][72],
reservoir_weight[58][73],
reservoir_weight[58][74],
reservoir_weight[58][75],
reservoir_weight[58][76],
reservoir_weight[58][77],
reservoir_weight[58][78],
reservoir_weight[58][79],
reservoir_weight[58][80],
reservoir_weight[58][81],
reservoir_weight[58][82],
reservoir_weight[58][83],
reservoir_weight[58][84],
reservoir_weight[58][85],
reservoir_weight[58][86],
reservoir_weight[58][87],
reservoir_weight[58][88],
reservoir_weight[58][89],
reservoir_weight[58][90],
reservoir_weight[58][91],
reservoir_weight[58][92],
reservoir_weight[58][93],
reservoir_weight[58][94],
reservoir_weight[58][95],
reservoir_weight[58][96],
reservoir_weight[58][97],
reservoir_weight[58][98],
reservoir_weight[58][99],
reservoir_weight[58][100],
reservoir_weight[58][101],
reservoir_weight[58][102],
reservoir_weight[58][103],
reservoir_weight[58][104],
reservoir_weight[58][105],
reservoir_weight[58][106],
reservoir_weight[58][107],
reservoir_weight[58][108],
reservoir_weight[58][109],
reservoir_weight[58][110],
reservoir_weight[58][111],
reservoir_weight[58][112],
reservoir_weight[58][113],
reservoir_weight[58][114],
reservoir_weight[58][115],
reservoir_weight[58][116],
reservoir_weight[58][117],
reservoir_weight[58][118],
reservoir_weight[58][119],
reservoir_weight[58][120],
reservoir_weight[58][121],
reservoir_weight[58][122],
reservoir_weight[58][123],
reservoir_weight[58][124],
reservoir_weight[58][125],
reservoir_weight[58][126],
reservoir_weight[58][127],
reservoir_weight[58][128],
reservoir_weight[58][129],
reservoir_weight[58][130],
reservoir_weight[58][131],
reservoir_weight[58][132],
reservoir_weight[58][133],
reservoir_weight[58][134],
reservoir_weight[58][135],
reservoir_weight[58][136],
reservoir_weight[58][137],
reservoir_weight[58][138],
reservoir_weight[58][139],
reservoir_weight[58][140],
reservoir_weight[58][141],
reservoir_weight[58][142],
reservoir_weight[58][143],
reservoir_weight[58][144],
reservoir_weight[58][145],
reservoir_weight[58][146],
reservoir_weight[58][147],
reservoir_weight[58][148],
reservoir_weight[58][149],
reservoir_weight[58][150],
reservoir_weight[58][151],
reservoir_weight[58][152],
reservoir_weight[58][153],
reservoir_weight[58][154],
reservoir_weight[58][155],
reservoir_weight[58][156],
reservoir_weight[58][157],
reservoir_weight[58][158],
reservoir_weight[58][159],
reservoir_weight[58][160],
reservoir_weight[58][161],
reservoir_weight[58][162],
reservoir_weight[58][163],
reservoir_weight[58][164],
reservoir_weight[58][165],
reservoir_weight[58][166],
reservoir_weight[58][167],
reservoir_weight[58][168],
reservoir_weight[58][169],
reservoir_weight[58][170],
reservoir_weight[58][171],
reservoir_weight[58][172],
reservoir_weight[58][173],
reservoir_weight[58][174],
reservoir_weight[58][175],
reservoir_weight[58][176],
reservoir_weight[58][177],
reservoir_weight[58][178],
reservoir_weight[58][179],
reservoir_weight[58][180],
reservoir_weight[58][181],
reservoir_weight[58][182],
reservoir_weight[58][183],
reservoir_weight[58][184],
reservoir_weight[58][185],
reservoir_weight[58][186],
reservoir_weight[58][187],
reservoir_weight[58][188],
reservoir_weight[58][189],
reservoir_weight[58][190],
reservoir_weight[58][191],
reservoir_weight[58][192],
reservoir_weight[58][193],
reservoir_weight[58][194],
reservoir_weight[58][195],
reservoir_weight[58][196],
reservoir_weight[58][197],
reservoir_weight[58][198],
reservoir_weight[58][199]
},
{reservoir_weight[59][0],
reservoir_weight[59][1],
reservoir_weight[59][2],
reservoir_weight[59][3],
reservoir_weight[59][4],
reservoir_weight[59][5],
reservoir_weight[59][6],
reservoir_weight[59][7],
reservoir_weight[59][8],
reservoir_weight[59][9],
reservoir_weight[59][10],
reservoir_weight[59][11],
reservoir_weight[59][12],
reservoir_weight[59][13],
reservoir_weight[59][14],
reservoir_weight[59][15],
reservoir_weight[59][16],
reservoir_weight[59][17],
reservoir_weight[59][18],
reservoir_weight[59][19],
reservoir_weight[59][20],
reservoir_weight[59][21],
reservoir_weight[59][22],
reservoir_weight[59][23],
reservoir_weight[59][24],
reservoir_weight[59][25],
reservoir_weight[59][26],
reservoir_weight[59][27],
reservoir_weight[59][28],
reservoir_weight[59][29],
reservoir_weight[59][30],
reservoir_weight[59][31],
reservoir_weight[59][32],
reservoir_weight[59][33],
reservoir_weight[59][34],
reservoir_weight[59][35],
reservoir_weight[59][36],
reservoir_weight[59][37],
reservoir_weight[59][38],
reservoir_weight[59][39],
reservoir_weight[59][40],
reservoir_weight[59][41],
reservoir_weight[59][42],
reservoir_weight[59][43],
reservoir_weight[59][44],
reservoir_weight[59][45],
reservoir_weight[59][46],
reservoir_weight[59][47],
reservoir_weight[59][48],
reservoir_weight[59][49],
reservoir_weight[59][50],
reservoir_weight[59][51],
reservoir_weight[59][52],
reservoir_weight[59][53],
reservoir_weight[59][54],
reservoir_weight[59][55],
reservoir_weight[59][56],
reservoir_weight[59][57],
reservoir_weight[59][58],
reservoir_weight[59][59],
reservoir_weight[59][60],
reservoir_weight[59][61],
reservoir_weight[59][62],
reservoir_weight[59][63],
reservoir_weight[59][64],
reservoir_weight[59][65],
reservoir_weight[59][66],
reservoir_weight[59][67],
reservoir_weight[59][68],
reservoir_weight[59][69],
reservoir_weight[59][70],
reservoir_weight[59][71],
reservoir_weight[59][72],
reservoir_weight[59][73],
reservoir_weight[59][74],
reservoir_weight[59][75],
reservoir_weight[59][76],
reservoir_weight[59][77],
reservoir_weight[59][78],
reservoir_weight[59][79],
reservoir_weight[59][80],
reservoir_weight[59][81],
reservoir_weight[59][82],
reservoir_weight[59][83],
reservoir_weight[59][84],
reservoir_weight[59][85],
reservoir_weight[59][86],
reservoir_weight[59][87],
reservoir_weight[59][88],
reservoir_weight[59][89],
reservoir_weight[59][90],
reservoir_weight[59][91],
reservoir_weight[59][92],
reservoir_weight[59][93],
reservoir_weight[59][94],
reservoir_weight[59][95],
reservoir_weight[59][96],
reservoir_weight[59][97],
reservoir_weight[59][98],
reservoir_weight[59][99],
reservoir_weight[59][100],
reservoir_weight[59][101],
reservoir_weight[59][102],
reservoir_weight[59][103],
reservoir_weight[59][104],
reservoir_weight[59][105],
reservoir_weight[59][106],
reservoir_weight[59][107],
reservoir_weight[59][108],
reservoir_weight[59][109],
reservoir_weight[59][110],
reservoir_weight[59][111],
reservoir_weight[59][112],
reservoir_weight[59][113],
reservoir_weight[59][114],
reservoir_weight[59][115],
reservoir_weight[59][116],
reservoir_weight[59][117],
reservoir_weight[59][118],
reservoir_weight[59][119],
reservoir_weight[59][120],
reservoir_weight[59][121],
reservoir_weight[59][122],
reservoir_weight[59][123],
reservoir_weight[59][124],
reservoir_weight[59][125],
reservoir_weight[59][126],
reservoir_weight[59][127],
reservoir_weight[59][128],
reservoir_weight[59][129],
reservoir_weight[59][130],
reservoir_weight[59][131],
reservoir_weight[59][132],
reservoir_weight[59][133],
reservoir_weight[59][134],
reservoir_weight[59][135],
reservoir_weight[59][136],
reservoir_weight[59][137],
reservoir_weight[59][138],
reservoir_weight[59][139],
reservoir_weight[59][140],
reservoir_weight[59][141],
reservoir_weight[59][142],
reservoir_weight[59][143],
reservoir_weight[59][144],
reservoir_weight[59][145],
reservoir_weight[59][146],
reservoir_weight[59][147],
reservoir_weight[59][148],
reservoir_weight[59][149],
reservoir_weight[59][150],
reservoir_weight[59][151],
reservoir_weight[59][152],
reservoir_weight[59][153],
reservoir_weight[59][154],
reservoir_weight[59][155],
reservoir_weight[59][156],
reservoir_weight[59][157],
reservoir_weight[59][158],
reservoir_weight[59][159],
reservoir_weight[59][160],
reservoir_weight[59][161],
reservoir_weight[59][162],
reservoir_weight[59][163],
reservoir_weight[59][164],
reservoir_weight[59][165],
reservoir_weight[59][166],
reservoir_weight[59][167],
reservoir_weight[59][168],
reservoir_weight[59][169],
reservoir_weight[59][170],
reservoir_weight[59][171],
reservoir_weight[59][172],
reservoir_weight[59][173],
reservoir_weight[59][174],
reservoir_weight[59][175],
reservoir_weight[59][176],
reservoir_weight[59][177],
reservoir_weight[59][178],
reservoir_weight[59][179],
reservoir_weight[59][180],
reservoir_weight[59][181],
reservoir_weight[59][182],
reservoir_weight[59][183],
reservoir_weight[59][184],
reservoir_weight[59][185],
reservoir_weight[59][186],
reservoir_weight[59][187],
reservoir_weight[59][188],
reservoir_weight[59][189],
reservoir_weight[59][190],
reservoir_weight[59][191],
reservoir_weight[59][192],
reservoir_weight[59][193],
reservoir_weight[59][194],
reservoir_weight[59][195],
reservoir_weight[59][196],
reservoir_weight[59][197],
reservoir_weight[59][198],
reservoir_weight[59][199]
},
{reservoir_weight[60][0],
reservoir_weight[60][1],
reservoir_weight[60][2],
reservoir_weight[60][3],
reservoir_weight[60][4],
reservoir_weight[60][5],
reservoir_weight[60][6],
reservoir_weight[60][7],
reservoir_weight[60][8],
reservoir_weight[60][9],
reservoir_weight[60][10],
reservoir_weight[60][11],
reservoir_weight[60][12],
reservoir_weight[60][13],
reservoir_weight[60][14],
reservoir_weight[60][15],
reservoir_weight[60][16],
reservoir_weight[60][17],
reservoir_weight[60][18],
reservoir_weight[60][19],
reservoir_weight[60][20],
reservoir_weight[60][21],
reservoir_weight[60][22],
reservoir_weight[60][23],
reservoir_weight[60][24],
reservoir_weight[60][25],
reservoir_weight[60][26],
reservoir_weight[60][27],
reservoir_weight[60][28],
reservoir_weight[60][29],
reservoir_weight[60][30],
reservoir_weight[60][31],
reservoir_weight[60][32],
reservoir_weight[60][33],
reservoir_weight[60][34],
reservoir_weight[60][35],
reservoir_weight[60][36],
reservoir_weight[60][37],
reservoir_weight[60][38],
reservoir_weight[60][39],
reservoir_weight[60][40],
reservoir_weight[60][41],
reservoir_weight[60][42],
reservoir_weight[60][43],
reservoir_weight[60][44],
reservoir_weight[60][45],
reservoir_weight[60][46],
reservoir_weight[60][47],
reservoir_weight[60][48],
reservoir_weight[60][49],
reservoir_weight[60][50],
reservoir_weight[60][51],
reservoir_weight[60][52],
reservoir_weight[60][53],
reservoir_weight[60][54],
reservoir_weight[60][55],
reservoir_weight[60][56],
reservoir_weight[60][57],
reservoir_weight[60][58],
reservoir_weight[60][59],
reservoir_weight[60][60],
reservoir_weight[60][61],
reservoir_weight[60][62],
reservoir_weight[60][63],
reservoir_weight[60][64],
reservoir_weight[60][65],
reservoir_weight[60][66],
reservoir_weight[60][67],
reservoir_weight[60][68],
reservoir_weight[60][69],
reservoir_weight[60][70],
reservoir_weight[60][71],
reservoir_weight[60][72],
reservoir_weight[60][73],
reservoir_weight[60][74],
reservoir_weight[60][75],
reservoir_weight[60][76],
reservoir_weight[60][77],
reservoir_weight[60][78],
reservoir_weight[60][79],
reservoir_weight[60][80],
reservoir_weight[60][81],
reservoir_weight[60][82],
reservoir_weight[60][83],
reservoir_weight[60][84],
reservoir_weight[60][85],
reservoir_weight[60][86],
reservoir_weight[60][87],
reservoir_weight[60][88],
reservoir_weight[60][89],
reservoir_weight[60][90],
reservoir_weight[60][91],
reservoir_weight[60][92],
reservoir_weight[60][93],
reservoir_weight[60][94],
reservoir_weight[60][95],
reservoir_weight[60][96],
reservoir_weight[60][97],
reservoir_weight[60][98],
reservoir_weight[60][99],
reservoir_weight[60][100],
reservoir_weight[60][101],
reservoir_weight[60][102],
reservoir_weight[60][103],
reservoir_weight[60][104],
reservoir_weight[60][105],
reservoir_weight[60][106],
reservoir_weight[60][107],
reservoir_weight[60][108],
reservoir_weight[60][109],
reservoir_weight[60][110],
reservoir_weight[60][111],
reservoir_weight[60][112],
reservoir_weight[60][113],
reservoir_weight[60][114],
reservoir_weight[60][115],
reservoir_weight[60][116],
reservoir_weight[60][117],
reservoir_weight[60][118],
reservoir_weight[60][119],
reservoir_weight[60][120],
reservoir_weight[60][121],
reservoir_weight[60][122],
reservoir_weight[60][123],
reservoir_weight[60][124],
reservoir_weight[60][125],
reservoir_weight[60][126],
reservoir_weight[60][127],
reservoir_weight[60][128],
reservoir_weight[60][129],
reservoir_weight[60][130],
reservoir_weight[60][131],
reservoir_weight[60][132],
reservoir_weight[60][133],
reservoir_weight[60][134],
reservoir_weight[60][135],
reservoir_weight[60][136],
reservoir_weight[60][137],
reservoir_weight[60][138],
reservoir_weight[60][139],
reservoir_weight[60][140],
reservoir_weight[60][141],
reservoir_weight[60][142],
reservoir_weight[60][143],
reservoir_weight[60][144],
reservoir_weight[60][145],
reservoir_weight[60][146],
reservoir_weight[60][147],
reservoir_weight[60][148],
reservoir_weight[60][149],
reservoir_weight[60][150],
reservoir_weight[60][151],
reservoir_weight[60][152],
reservoir_weight[60][153],
reservoir_weight[60][154],
reservoir_weight[60][155],
reservoir_weight[60][156],
reservoir_weight[60][157],
reservoir_weight[60][158],
reservoir_weight[60][159],
reservoir_weight[60][160],
reservoir_weight[60][161],
reservoir_weight[60][162],
reservoir_weight[60][163],
reservoir_weight[60][164],
reservoir_weight[60][165],
reservoir_weight[60][166],
reservoir_weight[60][167],
reservoir_weight[60][168],
reservoir_weight[60][169],
reservoir_weight[60][170],
reservoir_weight[60][171],
reservoir_weight[60][172],
reservoir_weight[60][173],
reservoir_weight[60][174],
reservoir_weight[60][175],
reservoir_weight[60][176],
reservoir_weight[60][177],
reservoir_weight[60][178],
reservoir_weight[60][179],
reservoir_weight[60][180],
reservoir_weight[60][181],
reservoir_weight[60][182],
reservoir_weight[60][183],
reservoir_weight[60][184],
reservoir_weight[60][185],
reservoir_weight[60][186],
reservoir_weight[60][187],
reservoir_weight[60][188],
reservoir_weight[60][189],
reservoir_weight[60][190],
reservoir_weight[60][191],
reservoir_weight[60][192],
reservoir_weight[60][193],
reservoir_weight[60][194],
reservoir_weight[60][195],
reservoir_weight[60][196],
reservoir_weight[60][197],
reservoir_weight[60][198],
reservoir_weight[60][199]
},
{reservoir_weight[61][0],
reservoir_weight[61][1],
reservoir_weight[61][2],
reservoir_weight[61][3],
reservoir_weight[61][4],
reservoir_weight[61][5],
reservoir_weight[61][6],
reservoir_weight[61][7],
reservoir_weight[61][8],
reservoir_weight[61][9],
reservoir_weight[61][10],
reservoir_weight[61][11],
reservoir_weight[61][12],
reservoir_weight[61][13],
reservoir_weight[61][14],
reservoir_weight[61][15],
reservoir_weight[61][16],
reservoir_weight[61][17],
reservoir_weight[61][18],
reservoir_weight[61][19],
reservoir_weight[61][20],
reservoir_weight[61][21],
reservoir_weight[61][22],
reservoir_weight[61][23],
reservoir_weight[61][24],
reservoir_weight[61][25],
reservoir_weight[61][26],
reservoir_weight[61][27],
reservoir_weight[61][28],
reservoir_weight[61][29],
reservoir_weight[61][30],
reservoir_weight[61][31],
reservoir_weight[61][32],
reservoir_weight[61][33],
reservoir_weight[61][34],
reservoir_weight[61][35],
reservoir_weight[61][36],
reservoir_weight[61][37],
reservoir_weight[61][38],
reservoir_weight[61][39],
reservoir_weight[61][40],
reservoir_weight[61][41],
reservoir_weight[61][42],
reservoir_weight[61][43],
reservoir_weight[61][44],
reservoir_weight[61][45],
reservoir_weight[61][46],
reservoir_weight[61][47],
reservoir_weight[61][48],
reservoir_weight[61][49],
reservoir_weight[61][50],
reservoir_weight[61][51],
reservoir_weight[61][52],
reservoir_weight[61][53],
reservoir_weight[61][54],
reservoir_weight[61][55],
reservoir_weight[61][56],
reservoir_weight[61][57],
reservoir_weight[61][58],
reservoir_weight[61][59],
reservoir_weight[61][60],
reservoir_weight[61][61],
reservoir_weight[61][62],
reservoir_weight[61][63],
reservoir_weight[61][64],
reservoir_weight[61][65],
reservoir_weight[61][66],
reservoir_weight[61][67],
reservoir_weight[61][68],
reservoir_weight[61][69],
reservoir_weight[61][70],
reservoir_weight[61][71],
reservoir_weight[61][72],
reservoir_weight[61][73],
reservoir_weight[61][74],
reservoir_weight[61][75],
reservoir_weight[61][76],
reservoir_weight[61][77],
reservoir_weight[61][78],
reservoir_weight[61][79],
reservoir_weight[61][80],
reservoir_weight[61][81],
reservoir_weight[61][82],
reservoir_weight[61][83],
reservoir_weight[61][84],
reservoir_weight[61][85],
reservoir_weight[61][86],
reservoir_weight[61][87],
reservoir_weight[61][88],
reservoir_weight[61][89],
reservoir_weight[61][90],
reservoir_weight[61][91],
reservoir_weight[61][92],
reservoir_weight[61][93],
reservoir_weight[61][94],
reservoir_weight[61][95],
reservoir_weight[61][96],
reservoir_weight[61][97],
reservoir_weight[61][98],
reservoir_weight[61][99],
reservoir_weight[61][100],
reservoir_weight[61][101],
reservoir_weight[61][102],
reservoir_weight[61][103],
reservoir_weight[61][104],
reservoir_weight[61][105],
reservoir_weight[61][106],
reservoir_weight[61][107],
reservoir_weight[61][108],
reservoir_weight[61][109],
reservoir_weight[61][110],
reservoir_weight[61][111],
reservoir_weight[61][112],
reservoir_weight[61][113],
reservoir_weight[61][114],
reservoir_weight[61][115],
reservoir_weight[61][116],
reservoir_weight[61][117],
reservoir_weight[61][118],
reservoir_weight[61][119],
reservoir_weight[61][120],
reservoir_weight[61][121],
reservoir_weight[61][122],
reservoir_weight[61][123],
reservoir_weight[61][124],
reservoir_weight[61][125],
reservoir_weight[61][126],
reservoir_weight[61][127],
reservoir_weight[61][128],
reservoir_weight[61][129],
reservoir_weight[61][130],
reservoir_weight[61][131],
reservoir_weight[61][132],
reservoir_weight[61][133],
reservoir_weight[61][134],
reservoir_weight[61][135],
reservoir_weight[61][136],
reservoir_weight[61][137],
reservoir_weight[61][138],
reservoir_weight[61][139],
reservoir_weight[61][140],
reservoir_weight[61][141],
reservoir_weight[61][142],
reservoir_weight[61][143],
reservoir_weight[61][144],
reservoir_weight[61][145],
reservoir_weight[61][146],
reservoir_weight[61][147],
reservoir_weight[61][148],
reservoir_weight[61][149],
reservoir_weight[61][150],
reservoir_weight[61][151],
reservoir_weight[61][152],
reservoir_weight[61][153],
reservoir_weight[61][154],
reservoir_weight[61][155],
reservoir_weight[61][156],
reservoir_weight[61][157],
reservoir_weight[61][158],
reservoir_weight[61][159],
reservoir_weight[61][160],
reservoir_weight[61][161],
reservoir_weight[61][162],
reservoir_weight[61][163],
reservoir_weight[61][164],
reservoir_weight[61][165],
reservoir_weight[61][166],
reservoir_weight[61][167],
reservoir_weight[61][168],
reservoir_weight[61][169],
reservoir_weight[61][170],
reservoir_weight[61][171],
reservoir_weight[61][172],
reservoir_weight[61][173],
reservoir_weight[61][174],
reservoir_weight[61][175],
reservoir_weight[61][176],
reservoir_weight[61][177],
reservoir_weight[61][178],
reservoir_weight[61][179],
reservoir_weight[61][180],
reservoir_weight[61][181],
reservoir_weight[61][182],
reservoir_weight[61][183],
reservoir_weight[61][184],
reservoir_weight[61][185],
reservoir_weight[61][186],
reservoir_weight[61][187],
reservoir_weight[61][188],
reservoir_weight[61][189],
reservoir_weight[61][190],
reservoir_weight[61][191],
reservoir_weight[61][192],
reservoir_weight[61][193],
reservoir_weight[61][194],
reservoir_weight[61][195],
reservoir_weight[61][196],
reservoir_weight[61][197],
reservoir_weight[61][198],
reservoir_weight[61][199]
},
{reservoir_weight[62][0],
reservoir_weight[62][1],
reservoir_weight[62][2],
reservoir_weight[62][3],
reservoir_weight[62][4],
reservoir_weight[62][5],
reservoir_weight[62][6],
reservoir_weight[62][7],
reservoir_weight[62][8],
reservoir_weight[62][9],
reservoir_weight[62][10],
reservoir_weight[62][11],
reservoir_weight[62][12],
reservoir_weight[62][13],
reservoir_weight[62][14],
reservoir_weight[62][15],
reservoir_weight[62][16],
reservoir_weight[62][17],
reservoir_weight[62][18],
reservoir_weight[62][19],
reservoir_weight[62][20],
reservoir_weight[62][21],
reservoir_weight[62][22],
reservoir_weight[62][23],
reservoir_weight[62][24],
reservoir_weight[62][25],
reservoir_weight[62][26],
reservoir_weight[62][27],
reservoir_weight[62][28],
reservoir_weight[62][29],
reservoir_weight[62][30],
reservoir_weight[62][31],
reservoir_weight[62][32],
reservoir_weight[62][33],
reservoir_weight[62][34],
reservoir_weight[62][35],
reservoir_weight[62][36],
reservoir_weight[62][37],
reservoir_weight[62][38],
reservoir_weight[62][39],
reservoir_weight[62][40],
reservoir_weight[62][41],
reservoir_weight[62][42],
reservoir_weight[62][43],
reservoir_weight[62][44],
reservoir_weight[62][45],
reservoir_weight[62][46],
reservoir_weight[62][47],
reservoir_weight[62][48],
reservoir_weight[62][49],
reservoir_weight[62][50],
reservoir_weight[62][51],
reservoir_weight[62][52],
reservoir_weight[62][53],
reservoir_weight[62][54],
reservoir_weight[62][55],
reservoir_weight[62][56],
reservoir_weight[62][57],
reservoir_weight[62][58],
reservoir_weight[62][59],
reservoir_weight[62][60],
reservoir_weight[62][61],
reservoir_weight[62][62],
reservoir_weight[62][63],
reservoir_weight[62][64],
reservoir_weight[62][65],
reservoir_weight[62][66],
reservoir_weight[62][67],
reservoir_weight[62][68],
reservoir_weight[62][69],
reservoir_weight[62][70],
reservoir_weight[62][71],
reservoir_weight[62][72],
reservoir_weight[62][73],
reservoir_weight[62][74],
reservoir_weight[62][75],
reservoir_weight[62][76],
reservoir_weight[62][77],
reservoir_weight[62][78],
reservoir_weight[62][79],
reservoir_weight[62][80],
reservoir_weight[62][81],
reservoir_weight[62][82],
reservoir_weight[62][83],
reservoir_weight[62][84],
reservoir_weight[62][85],
reservoir_weight[62][86],
reservoir_weight[62][87],
reservoir_weight[62][88],
reservoir_weight[62][89],
reservoir_weight[62][90],
reservoir_weight[62][91],
reservoir_weight[62][92],
reservoir_weight[62][93],
reservoir_weight[62][94],
reservoir_weight[62][95],
reservoir_weight[62][96],
reservoir_weight[62][97],
reservoir_weight[62][98],
reservoir_weight[62][99],
reservoir_weight[62][100],
reservoir_weight[62][101],
reservoir_weight[62][102],
reservoir_weight[62][103],
reservoir_weight[62][104],
reservoir_weight[62][105],
reservoir_weight[62][106],
reservoir_weight[62][107],
reservoir_weight[62][108],
reservoir_weight[62][109],
reservoir_weight[62][110],
reservoir_weight[62][111],
reservoir_weight[62][112],
reservoir_weight[62][113],
reservoir_weight[62][114],
reservoir_weight[62][115],
reservoir_weight[62][116],
reservoir_weight[62][117],
reservoir_weight[62][118],
reservoir_weight[62][119],
reservoir_weight[62][120],
reservoir_weight[62][121],
reservoir_weight[62][122],
reservoir_weight[62][123],
reservoir_weight[62][124],
reservoir_weight[62][125],
reservoir_weight[62][126],
reservoir_weight[62][127],
reservoir_weight[62][128],
reservoir_weight[62][129],
reservoir_weight[62][130],
reservoir_weight[62][131],
reservoir_weight[62][132],
reservoir_weight[62][133],
reservoir_weight[62][134],
reservoir_weight[62][135],
reservoir_weight[62][136],
reservoir_weight[62][137],
reservoir_weight[62][138],
reservoir_weight[62][139],
reservoir_weight[62][140],
reservoir_weight[62][141],
reservoir_weight[62][142],
reservoir_weight[62][143],
reservoir_weight[62][144],
reservoir_weight[62][145],
reservoir_weight[62][146],
reservoir_weight[62][147],
reservoir_weight[62][148],
reservoir_weight[62][149],
reservoir_weight[62][150],
reservoir_weight[62][151],
reservoir_weight[62][152],
reservoir_weight[62][153],
reservoir_weight[62][154],
reservoir_weight[62][155],
reservoir_weight[62][156],
reservoir_weight[62][157],
reservoir_weight[62][158],
reservoir_weight[62][159],
reservoir_weight[62][160],
reservoir_weight[62][161],
reservoir_weight[62][162],
reservoir_weight[62][163],
reservoir_weight[62][164],
reservoir_weight[62][165],
reservoir_weight[62][166],
reservoir_weight[62][167],
reservoir_weight[62][168],
reservoir_weight[62][169],
reservoir_weight[62][170],
reservoir_weight[62][171],
reservoir_weight[62][172],
reservoir_weight[62][173],
reservoir_weight[62][174],
reservoir_weight[62][175],
reservoir_weight[62][176],
reservoir_weight[62][177],
reservoir_weight[62][178],
reservoir_weight[62][179],
reservoir_weight[62][180],
reservoir_weight[62][181],
reservoir_weight[62][182],
reservoir_weight[62][183],
reservoir_weight[62][184],
reservoir_weight[62][185],
reservoir_weight[62][186],
reservoir_weight[62][187],
reservoir_weight[62][188],
reservoir_weight[62][189],
reservoir_weight[62][190],
reservoir_weight[62][191],
reservoir_weight[62][192],
reservoir_weight[62][193],
reservoir_weight[62][194],
reservoir_weight[62][195],
reservoir_weight[62][196],
reservoir_weight[62][197],
reservoir_weight[62][198],
reservoir_weight[62][199]
},
{reservoir_weight[63][0],
reservoir_weight[63][1],
reservoir_weight[63][2],
reservoir_weight[63][3],
reservoir_weight[63][4],
reservoir_weight[63][5],
reservoir_weight[63][6],
reservoir_weight[63][7],
reservoir_weight[63][8],
reservoir_weight[63][9],
reservoir_weight[63][10],
reservoir_weight[63][11],
reservoir_weight[63][12],
reservoir_weight[63][13],
reservoir_weight[63][14],
reservoir_weight[63][15],
reservoir_weight[63][16],
reservoir_weight[63][17],
reservoir_weight[63][18],
reservoir_weight[63][19],
reservoir_weight[63][20],
reservoir_weight[63][21],
reservoir_weight[63][22],
reservoir_weight[63][23],
reservoir_weight[63][24],
reservoir_weight[63][25],
reservoir_weight[63][26],
reservoir_weight[63][27],
reservoir_weight[63][28],
reservoir_weight[63][29],
reservoir_weight[63][30],
reservoir_weight[63][31],
reservoir_weight[63][32],
reservoir_weight[63][33],
reservoir_weight[63][34],
reservoir_weight[63][35],
reservoir_weight[63][36],
reservoir_weight[63][37],
reservoir_weight[63][38],
reservoir_weight[63][39],
reservoir_weight[63][40],
reservoir_weight[63][41],
reservoir_weight[63][42],
reservoir_weight[63][43],
reservoir_weight[63][44],
reservoir_weight[63][45],
reservoir_weight[63][46],
reservoir_weight[63][47],
reservoir_weight[63][48],
reservoir_weight[63][49],
reservoir_weight[63][50],
reservoir_weight[63][51],
reservoir_weight[63][52],
reservoir_weight[63][53],
reservoir_weight[63][54],
reservoir_weight[63][55],
reservoir_weight[63][56],
reservoir_weight[63][57],
reservoir_weight[63][58],
reservoir_weight[63][59],
reservoir_weight[63][60],
reservoir_weight[63][61],
reservoir_weight[63][62],
reservoir_weight[63][63],
reservoir_weight[63][64],
reservoir_weight[63][65],
reservoir_weight[63][66],
reservoir_weight[63][67],
reservoir_weight[63][68],
reservoir_weight[63][69],
reservoir_weight[63][70],
reservoir_weight[63][71],
reservoir_weight[63][72],
reservoir_weight[63][73],
reservoir_weight[63][74],
reservoir_weight[63][75],
reservoir_weight[63][76],
reservoir_weight[63][77],
reservoir_weight[63][78],
reservoir_weight[63][79],
reservoir_weight[63][80],
reservoir_weight[63][81],
reservoir_weight[63][82],
reservoir_weight[63][83],
reservoir_weight[63][84],
reservoir_weight[63][85],
reservoir_weight[63][86],
reservoir_weight[63][87],
reservoir_weight[63][88],
reservoir_weight[63][89],
reservoir_weight[63][90],
reservoir_weight[63][91],
reservoir_weight[63][92],
reservoir_weight[63][93],
reservoir_weight[63][94],
reservoir_weight[63][95],
reservoir_weight[63][96],
reservoir_weight[63][97],
reservoir_weight[63][98],
reservoir_weight[63][99],
reservoir_weight[63][100],
reservoir_weight[63][101],
reservoir_weight[63][102],
reservoir_weight[63][103],
reservoir_weight[63][104],
reservoir_weight[63][105],
reservoir_weight[63][106],
reservoir_weight[63][107],
reservoir_weight[63][108],
reservoir_weight[63][109],
reservoir_weight[63][110],
reservoir_weight[63][111],
reservoir_weight[63][112],
reservoir_weight[63][113],
reservoir_weight[63][114],
reservoir_weight[63][115],
reservoir_weight[63][116],
reservoir_weight[63][117],
reservoir_weight[63][118],
reservoir_weight[63][119],
reservoir_weight[63][120],
reservoir_weight[63][121],
reservoir_weight[63][122],
reservoir_weight[63][123],
reservoir_weight[63][124],
reservoir_weight[63][125],
reservoir_weight[63][126],
reservoir_weight[63][127],
reservoir_weight[63][128],
reservoir_weight[63][129],
reservoir_weight[63][130],
reservoir_weight[63][131],
reservoir_weight[63][132],
reservoir_weight[63][133],
reservoir_weight[63][134],
reservoir_weight[63][135],
reservoir_weight[63][136],
reservoir_weight[63][137],
reservoir_weight[63][138],
reservoir_weight[63][139],
reservoir_weight[63][140],
reservoir_weight[63][141],
reservoir_weight[63][142],
reservoir_weight[63][143],
reservoir_weight[63][144],
reservoir_weight[63][145],
reservoir_weight[63][146],
reservoir_weight[63][147],
reservoir_weight[63][148],
reservoir_weight[63][149],
reservoir_weight[63][150],
reservoir_weight[63][151],
reservoir_weight[63][152],
reservoir_weight[63][153],
reservoir_weight[63][154],
reservoir_weight[63][155],
reservoir_weight[63][156],
reservoir_weight[63][157],
reservoir_weight[63][158],
reservoir_weight[63][159],
reservoir_weight[63][160],
reservoir_weight[63][161],
reservoir_weight[63][162],
reservoir_weight[63][163],
reservoir_weight[63][164],
reservoir_weight[63][165],
reservoir_weight[63][166],
reservoir_weight[63][167],
reservoir_weight[63][168],
reservoir_weight[63][169],
reservoir_weight[63][170],
reservoir_weight[63][171],
reservoir_weight[63][172],
reservoir_weight[63][173],
reservoir_weight[63][174],
reservoir_weight[63][175],
reservoir_weight[63][176],
reservoir_weight[63][177],
reservoir_weight[63][178],
reservoir_weight[63][179],
reservoir_weight[63][180],
reservoir_weight[63][181],
reservoir_weight[63][182],
reservoir_weight[63][183],
reservoir_weight[63][184],
reservoir_weight[63][185],
reservoir_weight[63][186],
reservoir_weight[63][187],
reservoir_weight[63][188],
reservoir_weight[63][189],
reservoir_weight[63][190],
reservoir_weight[63][191],
reservoir_weight[63][192],
reservoir_weight[63][193],
reservoir_weight[63][194],
reservoir_weight[63][195],
reservoir_weight[63][196],
reservoir_weight[63][197],
reservoir_weight[63][198],
reservoir_weight[63][199]
},
{reservoir_weight[64][0],
reservoir_weight[64][1],
reservoir_weight[64][2],
reservoir_weight[64][3],
reservoir_weight[64][4],
reservoir_weight[64][5],
reservoir_weight[64][6],
reservoir_weight[64][7],
reservoir_weight[64][8],
reservoir_weight[64][9],
reservoir_weight[64][10],
reservoir_weight[64][11],
reservoir_weight[64][12],
reservoir_weight[64][13],
reservoir_weight[64][14],
reservoir_weight[64][15],
reservoir_weight[64][16],
reservoir_weight[64][17],
reservoir_weight[64][18],
reservoir_weight[64][19],
reservoir_weight[64][20],
reservoir_weight[64][21],
reservoir_weight[64][22],
reservoir_weight[64][23],
reservoir_weight[64][24],
reservoir_weight[64][25],
reservoir_weight[64][26],
reservoir_weight[64][27],
reservoir_weight[64][28],
reservoir_weight[64][29],
reservoir_weight[64][30],
reservoir_weight[64][31],
reservoir_weight[64][32],
reservoir_weight[64][33],
reservoir_weight[64][34],
reservoir_weight[64][35],
reservoir_weight[64][36],
reservoir_weight[64][37],
reservoir_weight[64][38],
reservoir_weight[64][39],
reservoir_weight[64][40],
reservoir_weight[64][41],
reservoir_weight[64][42],
reservoir_weight[64][43],
reservoir_weight[64][44],
reservoir_weight[64][45],
reservoir_weight[64][46],
reservoir_weight[64][47],
reservoir_weight[64][48],
reservoir_weight[64][49],
reservoir_weight[64][50],
reservoir_weight[64][51],
reservoir_weight[64][52],
reservoir_weight[64][53],
reservoir_weight[64][54],
reservoir_weight[64][55],
reservoir_weight[64][56],
reservoir_weight[64][57],
reservoir_weight[64][58],
reservoir_weight[64][59],
reservoir_weight[64][60],
reservoir_weight[64][61],
reservoir_weight[64][62],
reservoir_weight[64][63],
reservoir_weight[64][64],
reservoir_weight[64][65],
reservoir_weight[64][66],
reservoir_weight[64][67],
reservoir_weight[64][68],
reservoir_weight[64][69],
reservoir_weight[64][70],
reservoir_weight[64][71],
reservoir_weight[64][72],
reservoir_weight[64][73],
reservoir_weight[64][74],
reservoir_weight[64][75],
reservoir_weight[64][76],
reservoir_weight[64][77],
reservoir_weight[64][78],
reservoir_weight[64][79],
reservoir_weight[64][80],
reservoir_weight[64][81],
reservoir_weight[64][82],
reservoir_weight[64][83],
reservoir_weight[64][84],
reservoir_weight[64][85],
reservoir_weight[64][86],
reservoir_weight[64][87],
reservoir_weight[64][88],
reservoir_weight[64][89],
reservoir_weight[64][90],
reservoir_weight[64][91],
reservoir_weight[64][92],
reservoir_weight[64][93],
reservoir_weight[64][94],
reservoir_weight[64][95],
reservoir_weight[64][96],
reservoir_weight[64][97],
reservoir_weight[64][98],
reservoir_weight[64][99],
reservoir_weight[64][100],
reservoir_weight[64][101],
reservoir_weight[64][102],
reservoir_weight[64][103],
reservoir_weight[64][104],
reservoir_weight[64][105],
reservoir_weight[64][106],
reservoir_weight[64][107],
reservoir_weight[64][108],
reservoir_weight[64][109],
reservoir_weight[64][110],
reservoir_weight[64][111],
reservoir_weight[64][112],
reservoir_weight[64][113],
reservoir_weight[64][114],
reservoir_weight[64][115],
reservoir_weight[64][116],
reservoir_weight[64][117],
reservoir_weight[64][118],
reservoir_weight[64][119],
reservoir_weight[64][120],
reservoir_weight[64][121],
reservoir_weight[64][122],
reservoir_weight[64][123],
reservoir_weight[64][124],
reservoir_weight[64][125],
reservoir_weight[64][126],
reservoir_weight[64][127],
reservoir_weight[64][128],
reservoir_weight[64][129],
reservoir_weight[64][130],
reservoir_weight[64][131],
reservoir_weight[64][132],
reservoir_weight[64][133],
reservoir_weight[64][134],
reservoir_weight[64][135],
reservoir_weight[64][136],
reservoir_weight[64][137],
reservoir_weight[64][138],
reservoir_weight[64][139],
reservoir_weight[64][140],
reservoir_weight[64][141],
reservoir_weight[64][142],
reservoir_weight[64][143],
reservoir_weight[64][144],
reservoir_weight[64][145],
reservoir_weight[64][146],
reservoir_weight[64][147],
reservoir_weight[64][148],
reservoir_weight[64][149],
reservoir_weight[64][150],
reservoir_weight[64][151],
reservoir_weight[64][152],
reservoir_weight[64][153],
reservoir_weight[64][154],
reservoir_weight[64][155],
reservoir_weight[64][156],
reservoir_weight[64][157],
reservoir_weight[64][158],
reservoir_weight[64][159],
reservoir_weight[64][160],
reservoir_weight[64][161],
reservoir_weight[64][162],
reservoir_weight[64][163],
reservoir_weight[64][164],
reservoir_weight[64][165],
reservoir_weight[64][166],
reservoir_weight[64][167],
reservoir_weight[64][168],
reservoir_weight[64][169],
reservoir_weight[64][170],
reservoir_weight[64][171],
reservoir_weight[64][172],
reservoir_weight[64][173],
reservoir_weight[64][174],
reservoir_weight[64][175],
reservoir_weight[64][176],
reservoir_weight[64][177],
reservoir_weight[64][178],
reservoir_weight[64][179],
reservoir_weight[64][180],
reservoir_weight[64][181],
reservoir_weight[64][182],
reservoir_weight[64][183],
reservoir_weight[64][184],
reservoir_weight[64][185],
reservoir_weight[64][186],
reservoir_weight[64][187],
reservoir_weight[64][188],
reservoir_weight[64][189],
reservoir_weight[64][190],
reservoir_weight[64][191],
reservoir_weight[64][192],
reservoir_weight[64][193],
reservoir_weight[64][194],
reservoir_weight[64][195],
reservoir_weight[64][196],
reservoir_weight[64][197],
reservoir_weight[64][198],
reservoir_weight[64][199]
},
{reservoir_weight[65][0],
reservoir_weight[65][1],
reservoir_weight[65][2],
reservoir_weight[65][3],
reservoir_weight[65][4],
reservoir_weight[65][5],
reservoir_weight[65][6],
reservoir_weight[65][7],
reservoir_weight[65][8],
reservoir_weight[65][9],
reservoir_weight[65][10],
reservoir_weight[65][11],
reservoir_weight[65][12],
reservoir_weight[65][13],
reservoir_weight[65][14],
reservoir_weight[65][15],
reservoir_weight[65][16],
reservoir_weight[65][17],
reservoir_weight[65][18],
reservoir_weight[65][19],
reservoir_weight[65][20],
reservoir_weight[65][21],
reservoir_weight[65][22],
reservoir_weight[65][23],
reservoir_weight[65][24],
reservoir_weight[65][25],
reservoir_weight[65][26],
reservoir_weight[65][27],
reservoir_weight[65][28],
reservoir_weight[65][29],
reservoir_weight[65][30],
reservoir_weight[65][31],
reservoir_weight[65][32],
reservoir_weight[65][33],
reservoir_weight[65][34],
reservoir_weight[65][35],
reservoir_weight[65][36],
reservoir_weight[65][37],
reservoir_weight[65][38],
reservoir_weight[65][39],
reservoir_weight[65][40],
reservoir_weight[65][41],
reservoir_weight[65][42],
reservoir_weight[65][43],
reservoir_weight[65][44],
reservoir_weight[65][45],
reservoir_weight[65][46],
reservoir_weight[65][47],
reservoir_weight[65][48],
reservoir_weight[65][49],
reservoir_weight[65][50],
reservoir_weight[65][51],
reservoir_weight[65][52],
reservoir_weight[65][53],
reservoir_weight[65][54],
reservoir_weight[65][55],
reservoir_weight[65][56],
reservoir_weight[65][57],
reservoir_weight[65][58],
reservoir_weight[65][59],
reservoir_weight[65][60],
reservoir_weight[65][61],
reservoir_weight[65][62],
reservoir_weight[65][63],
reservoir_weight[65][64],
reservoir_weight[65][65],
reservoir_weight[65][66],
reservoir_weight[65][67],
reservoir_weight[65][68],
reservoir_weight[65][69],
reservoir_weight[65][70],
reservoir_weight[65][71],
reservoir_weight[65][72],
reservoir_weight[65][73],
reservoir_weight[65][74],
reservoir_weight[65][75],
reservoir_weight[65][76],
reservoir_weight[65][77],
reservoir_weight[65][78],
reservoir_weight[65][79],
reservoir_weight[65][80],
reservoir_weight[65][81],
reservoir_weight[65][82],
reservoir_weight[65][83],
reservoir_weight[65][84],
reservoir_weight[65][85],
reservoir_weight[65][86],
reservoir_weight[65][87],
reservoir_weight[65][88],
reservoir_weight[65][89],
reservoir_weight[65][90],
reservoir_weight[65][91],
reservoir_weight[65][92],
reservoir_weight[65][93],
reservoir_weight[65][94],
reservoir_weight[65][95],
reservoir_weight[65][96],
reservoir_weight[65][97],
reservoir_weight[65][98],
reservoir_weight[65][99],
reservoir_weight[65][100],
reservoir_weight[65][101],
reservoir_weight[65][102],
reservoir_weight[65][103],
reservoir_weight[65][104],
reservoir_weight[65][105],
reservoir_weight[65][106],
reservoir_weight[65][107],
reservoir_weight[65][108],
reservoir_weight[65][109],
reservoir_weight[65][110],
reservoir_weight[65][111],
reservoir_weight[65][112],
reservoir_weight[65][113],
reservoir_weight[65][114],
reservoir_weight[65][115],
reservoir_weight[65][116],
reservoir_weight[65][117],
reservoir_weight[65][118],
reservoir_weight[65][119],
reservoir_weight[65][120],
reservoir_weight[65][121],
reservoir_weight[65][122],
reservoir_weight[65][123],
reservoir_weight[65][124],
reservoir_weight[65][125],
reservoir_weight[65][126],
reservoir_weight[65][127],
reservoir_weight[65][128],
reservoir_weight[65][129],
reservoir_weight[65][130],
reservoir_weight[65][131],
reservoir_weight[65][132],
reservoir_weight[65][133],
reservoir_weight[65][134],
reservoir_weight[65][135],
reservoir_weight[65][136],
reservoir_weight[65][137],
reservoir_weight[65][138],
reservoir_weight[65][139],
reservoir_weight[65][140],
reservoir_weight[65][141],
reservoir_weight[65][142],
reservoir_weight[65][143],
reservoir_weight[65][144],
reservoir_weight[65][145],
reservoir_weight[65][146],
reservoir_weight[65][147],
reservoir_weight[65][148],
reservoir_weight[65][149],
reservoir_weight[65][150],
reservoir_weight[65][151],
reservoir_weight[65][152],
reservoir_weight[65][153],
reservoir_weight[65][154],
reservoir_weight[65][155],
reservoir_weight[65][156],
reservoir_weight[65][157],
reservoir_weight[65][158],
reservoir_weight[65][159],
reservoir_weight[65][160],
reservoir_weight[65][161],
reservoir_weight[65][162],
reservoir_weight[65][163],
reservoir_weight[65][164],
reservoir_weight[65][165],
reservoir_weight[65][166],
reservoir_weight[65][167],
reservoir_weight[65][168],
reservoir_weight[65][169],
reservoir_weight[65][170],
reservoir_weight[65][171],
reservoir_weight[65][172],
reservoir_weight[65][173],
reservoir_weight[65][174],
reservoir_weight[65][175],
reservoir_weight[65][176],
reservoir_weight[65][177],
reservoir_weight[65][178],
reservoir_weight[65][179],
reservoir_weight[65][180],
reservoir_weight[65][181],
reservoir_weight[65][182],
reservoir_weight[65][183],
reservoir_weight[65][184],
reservoir_weight[65][185],
reservoir_weight[65][186],
reservoir_weight[65][187],
reservoir_weight[65][188],
reservoir_weight[65][189],
reservoir_weight[65][190],
reservoir_weight[65][191],
reservoir_weight[65][192],
reservoir_weight[65][193],
reservoir_weight[65][194],
reservoir_weight[65][195],
reservoir_weight[65][196],
reservoir_weight[65][197],
reservoir_weight[65][198],
reservoir_weight[65][199]
},
{reservoir_weight[66][0],
reservoir_weight[66][1],
reservoir_weight[66][2],
reservoir_weight[66][3],
reservoir_weight[66][4],
reservoir_weight[66][5],
reservoir_weight[66][6],
reservoir_weight[66][7],
reservoir_weight[66][8],
reservoir_weight[66][9],
reservoir_weight[66][10],
reservoir_weight[66][11],
reservoir_weight[66][12],
reservoir_weight[66][13],
reservoir_weight[66][14],
reservoir_weight[66][15],
reservoir_weight[66][16],
reservoir_weight[66][17],
reservoir_weight[66][18],
reservoir_weight[66][19],
reservoir_weight[66][20],
reservoir_weight[66][21],
reservoir_weight[66][22],
reservoir_weight[66][23],
reservoir_weight[66][24],
reservoir_weight[66][25],
reservoir_weight[66][26],
reservoir_weight[66][27],
reservoir_weight[66][28],
reservoir_weight[66][29],
reservoir_weight[66][30],
reservoir_weight[66][31],
reservoir_weight[66][32],
reservoir_weight[66][33],
reservoir_weight[66][34],
reservoir_weight[66][35],
reservoir_weight[66][36],
reservoir_weight[66][37],
reservoir_weight[66][38],
reservoir_weight[66][39],
reservoir_weight[66][40],
reservoir_weight[66][41],
reservoir_weight[66][42],
reservoir_weight[66][43],
reservoir_weight[66][44],
reservoir_weight[66][45],
reservoir_weight[66][46],
reservoir_weight[66][47],
reservoir_weight[66][48],
reservoir_weight[66][49],
reservoir_weight[66][50],
reservoir_weight[66][51],
reservoir_weight[66][52],
reservoir_weight[66][53],
reservoir_weight[66][54],
reservoir_weight[66][55],
reservoir_weight[66][56],
reservoir_weight[66][57],
reservoir_weight[66][58],
reservoir_weight[66][59],
reservoir_weight[66][60],
reservoir_weight[66][61],
reservoir_weight[66][62],
reservoir_weight[66][63],
reservoir_weight[66][64],
reservoir_weight[66][65],
reservoir_weight[66][66],
reservoir_weight[66][67],
reservoir_weight[66][68],
reservoir_weight[66][69],
reservoir_weight[66][70],
reservoir_weight[66][71],
reservoir_weight[66][72],
reservoir_weight[66][73],
reservoir_weight[66][74],
reservoir_weight[66][75],
reservoir_weight[66][76],
reservoir_weight[66][77],
reservoir_weight[66][78],
reservoir_weight[66][79],
reservoir_weight[66][80],
reservoir_weight[66][81],
reservoir_weight[66][82],
reservoir_weight[66][83],
reservoir_weight[66][84],
reservoir_weight[66][85],
reservoir_weight[66][86],
reservoir_weight[66][87],
reservoir_weight[66][88],
reservoir_weight[66][89],
reservoir_weight[66][90],
reservoir_weight[66][91],
reservoir_weight[66][92],
reservoir_weight[66][93],
reservoir_weight[66][94],
reservoir_weight[66][95],
reservoir_weight[66][96],
reservoir_weight[66][97],
reservoir_weight[66][98],
reservoir_weight[66][99],
reservoir_weight[66][100],
reservoir_weight[66][101],
reservoir_weight[66][102],
reservoir_weight[66][103],
reservoir_weight[66][104],
reservoir_weight[66][105],
reservoir_weight[66][106],
reservoir_weight[66][107],
reservoir_weight[66][108],
reservoir_weight[66][109],
reservoir_weight[66][110],
reservoir_weight[66][111],
reservoir_weight[66][112],
reservoir_weight[66][113],
reservoir_weight[66][114],
reservoir_weight[66][115],
reservoir_weight[66][116],
reservoir_weight[66][117],
reservoir_weight[66][118],
reservoir_weight[66][119],
reservoir_weight[66][120],
reservoir_weight[66][121],
reservoir_weight[66][122],
reservoir_weight[66][123],
reservoir_weight[66][124],
reservoir_weight[66][125],
reservoir_weight[66][126],
reservoir_weight[66][127],
reservoir_weight[66][128],
reservoir_weight[66][129],
reservoir_weight[66][130],
reservoir_weight[66][131],
reservoir_weight[66][132],
reservoir_weight[66][133],
reservoir_weight[66][134],
reservoir_weight[66][135],
reservoir_weight[66][136],
reservoir_weight[66][137],
reservoir_weight[66][138],
reservoir_weight[66][139],
reservoir_weight[66][140],
reservoir_weight[66][141],
reservoir_weight[66][142],
reservoir_weight[66][143],
reservoir_weight[66][144],
reservoir_weight[66][145],
reservoir_weight[66][146],
reservoir_weight[66][147],
reservoir_weight[66][148],
reservoir_weight[66][149],
reservoir_weight[66][150],
reservoir_weight[66][151],
reservoir_weight[66][152],
reservoir_weight[66][153],
reservoir_weight[66][154],
reservoir_weight[66][155],
reservoir_weight[66][156],
reservoir_weight[66][157],
reservoir_weight[66][158],
reservoir_weight[66][159],
reservoir_weight[66][160],
reservoir_weight[66][161],
reservoir_weight[66][162],
reservoir_weight[66][163],
reservoir_weight[66][164],
reservoir_weight[66][165],
reservoir_weight[66][166],
reservoir_weight[66][167],
reservoir_weight[66][168],
reservoir_weight[66][169],
reservoir_weight[66][170],
reservoir_weight[66][171],
reservoir_weight[66][172],
reservoir_weight[66][173],
reservoir_weight[66][174],
reservoir_weight[66][175],
reservoir_weight[66][176],
reservoir_weight[66][177],
reservoir_weight[66][178],
reservoir_weight[66][179],
reservoir_weight[66][180],
reservoir_weight[66][181],
reservoir_weight[66][182],
reservoir_weight[66][183],
reservoir_weight[66][184],
reservoir_weight[66][185],
reservoir_weight[66][186],
reservoir_weight[66][187],
reservoir_weight[66][188],
reservoir_weight[66][189],
reservoir_weight[66][190],
reservoir_weight[66][191],
reservoir_weight[66][192],
reservoir_weight[66][193],
reservoir_weight[66][194],
reservoir_weight[66][195],
reservoir_weight[66][196],
reservoir_weight[66][197],
reservoir_weight[66][198],
reservoir_weight[66][199]
},
{reservoir_weight[67][0],
reservoir_weight[67][1],
reservoir_weight[67][2],
reservoir_weight[67][3],
reservoir_weight[67][4],
reservoir_weight[67][5],
reservoir_weight[67][6],
reservoir_weight[67][7],
reservoir_weight[67][8],
reservoir_weight[67][9],
reservoir_weight[67][10],
reservoir_weight[67][11],
reservoir_weight[67][12],
reservoir_weight[67][13],
reservoir_weight[67][14],
reservoir_weight[67][15],
reservoir_weight[67][16],
reservoir_weight[67][17],
reservoir_weight[67][18],
reservoir_weight[67][19],
reservoir_weight[67][20],
reservoir_weight[67][21],
reservoir_weight[67][22],
reservoir_weight[67][23],
reservoir_weight[67][24],
reservoir_weight[67][25],
reservoir_weight[67][26],
reservoir_weight[67][27],
reservoir_weight[67][28],
reservoir_weight[67][29],
reservoir_weight[67][30],
reservoir_weight[67][31],
reservoir_weight[67][32],
reservoir_weight[67][33],
reservoir_weight[67][34],
reservoir_weight[67][35],
reservoir_weight[67][36],
reservoir_weight[67][37],
reservoir_weight[67][38],
reservoir_weight[67][39],
reservoir_weight[67][40],
reservoir_weight[67][41],
reservoir_weight[67][42],
reservoir_weight[67][43],
reservoir_weight[67][44],
reservoir_weight[67][45],
reservoir_weight[67][46],
reservoir_weight[67][47],
reservoir_weight[67][48],
reservoir_weight[67][49],
reservoir_weight[67][50],
reservoir_weight[67][51],
reservoir_weight[67][52],
reservoir_weight[67][53],
reservoir_weight[67][54],
reservoir_weight[67][55],
reservoir_weight[67][56],
reservoir_weight[67][57],
reservoir_weight[67][58],
reservoir_weight[67][59],
reservoir_weight[67][60],
reservoir_weight[67][61],
reservoir_weight[67][62],
reservoir_weight[67][63],
reservoir_weight[67][64],
reservoir_weight[67][65],
reservoir_weight[67][66],
reservoir_weight[67][67],
reservoir_weight[67][68],
reservoir_weight[67][69],
reservoir_weight[67][70],
reservoir_weight[67][71],
reservoir_weight[67][72],
reservoir_weight[67][73],
reservoir_weight[67][74],
reservoir_weight[67][75],
reservoir_weight[67][76],
reservoir_weight[67][77],
reservoir_weight[67][78],
reservoir_weight[67][79],
reservoir_weight[67][80],
reservoir_weight[67][81],
reservoir_weight[67][82],
reservoir_weight[67][83],
reservoir_weight[67][84],
reservoir_weight[67][85],
reservoir_weight[67][86],
reservoir_weight[67][87],
reservoir_weight[67][88],
reservoir_weight[67][89],
reservoir_weight[67][90],
reservoir_weight[67][91],
reservoir_weight[67][92],
reservoir_weight[67][93],
reservoir_weight[67][94],
reservoir_weight[67][95],
reservoir_weight[67][96],
reservoir_weight[67][97],
reservoir_weight[67][98],
reservoir_weight[67][99],
reservoir_weight[67][100],
reservoir_weight[67][101],
reservoir_weight[67][102],
reservoir_weight[67][103],
reservoir_weight[67][104],
reservoir_weight[67][105],
reservoir_weight[67][106],
reservoir_weight[67][107],
reservoir_weight[67][108],
reservoir_weight[67][109],
reservoir_weight[67][110],
reservoir_weight[67][111],
reservoir_weight[67][112],
reservoir_weight[67][113],
reservoir_weight[67][114],
reservoir_weight[67][115],
reservoir_weight[67][116],
reservoir_weight[67][117],
reservoir_weight[67][118],
reservoir_weight[67][119],
reservoir_weight[67][120],
reservoir_weight[67][121],
reservoir_weight[67][122],
reservoir_weight[67][123],
reservoir_weight[67][124],
reservoir_weight[67][125],
reservoir_weight[67][126],
reservoir_weight[67][127],
reservoir_weight[67][128],
reservoir_weight[67][129],
reservoir_weight[67][130],
reservoir_weight[67][131],
reservoir_weight[67][132],
reservoir_weight[67][133],
reservoir_weight[67][134],
reservoir_weight[67][135],
reservoir_weight[67][136],
reservoir_weight[67][137],
reservoir_weight[67][138],
reservoir_weight[67][139],
reservoir_weight[67][140],
reservoir_weight[67][141],
reservoir_weight[67][142],
reservoir_weight[67][143],
reservoir_weight[67][144],
reservoir_weight[67][145],
reservoir_weight[67][146],
reservoir_weight[67][147],
reservoir_weight[67][148],
reservoir_weight[67][149],
reservoir_weight[67][150],
reservoir_weight[67][151],
reservoir_weight[67][152],
reservoir_weight[67][153],
reservoir_weight[67][154],
reservoir_weight[67][155],
reservoir_weight[67][156],
reservoir_weight[67][157],
reservoir_weight[67][158],
reservoir_weight[67][159],
reservoir_weight[67][160],
reservoir_weight[67][161],
reservoir_weight[67][162],
reservoir_weight[67][163],
reservoir_weight[67][164],
reservoir_weight[67][165],
reservoir_weight[67][166],
reservoir_weight[67][167],
reservoir_weight[67][168],
reservoir_weight[67][169],
reservoir_weight[67][170],
reservoir_weight[67][171],
reservoir_weight[67][172],
reservoir_weight[67][173],
reservoir_weight[67][174],
reservoir_weight[67][175],
reservoir_weight[67][176],
reservoir_weight[67][177],
reservoir_weight[67][178],
reservoir_weight[67][179],
reservoir_weight[67][180],
reservoir_weight[67][181],
reservoir_weight[67][182],
reservoir_weight[67][183],
reservoir_weight[67][184],
reservoir_weight[67][185],
reservoir_weight[67][186],
reservoir_weight[67][187],
reservoir_weight[67][188],
reservoir_weight[67][189],
reservoir_weight[67][190],
reservoir_weight[67][191],
reservoir_weight[67][192],
reservoir_weight[67][193],
reservoir_weight[67][194],
reservoir_weight[67][195],
reservoir_weight[67][196],
reservoir_weight[67][197],
reservoir_weight[67][198],
reservoir_weight[67][199]
},
{reservoir_weight[68][0],
reservoir_weight[68][1],
reservoir_weight[68][2],
reservoir_weight[68][3],
reservoir_weight[68][4],
reservoir_weight[68][5],
reservoir_weight[68][6],
reservoir_weight[68][7],
reservoir_weight[68][8],
reservoir_weight[68][9],
reservoir_weight[68][10],
reservoir_weight[68][11],
reservoir_weight[68][12],
reservoir_weight[68][13],
reservoir_weight[68][14],
reservoir_weight[68][15],
reservoir_weight[68][16],
reservoir_weight[68][17],
reservoir_weight[68][18],
reservoir_weight[68][19],
reservoir_weight[68][20],
reservoir_weight[68][21],
reservoir_weight[68][22],
reservoir_weight[68][23],
reservoir_weight[68][24],
reservoir_weight[68][25],
reservoir_weight[68][26],
reservoir_weight[68][27],
reservoir_weight[68][28],
reservoir_weight[68][29],
reservoir_weight[68][30],
reservoir_weight[68][31],
reservoir_weight[68][32],
reservoir_weight[68][33],
reservoir_weight[68][34],
reservoir_weight[68][35],
reservoir_weight[68][36],
reservoir_weight[68][37],
reservoir_weight[68][38],
reservoir_weight[68][39],
reservoir_weight[68][40],
reservoir_weight[68][41],
reservoir_weight[68][42],
reservoir_weight[68][43],
reservoir_weight[68][44],
reservoir_weight[68][45],
reservoir_weight[68][46],
reservoir_weight[68][47],
reservoir_weight[68][48],
reservoir_weight[68][49],
reservoir_weight[68][50],
reservoir_weight[68][51],
reservoir_weight[68][52],
reservoir_weight[68][53],
reservoir_weight[68][54],
reservoir_weight[68][55],
reservoir_weight[68][56],
reservoir_weight[68][57],
reservoir_weight[68][58],
reservoir_weight[68][59],
reservoir_weight[68][60],
reservoir_weight[68][61],
reservoir_weight[68][62],
reservoir_weight[68][63],
reservoir_weight[68][64],
reservoir_weight[68][65],
reservoir_weight[68][66],
reservoir_weight[68][67],
reservoir_weight[68][68],
reservoir_weight[68][69],
reservoir_weight[68][70],
reservoir_weight[68][71],
reservoir_weight[68][72],
reservoir_weight[68][73],
reservoir_weight[68][74],
reservoir_weight[68][75],
reservoir_weight[68][76],
reservoir_weight[68][77],
reservoir_weight[68][78],
reservoir_weight[68][79],
reservoir_weight[68][80],
reservoir_weight[68][81],
reservoir_weight[68][82],
reservoir_weight[68][83],
reservoir_weight[68][84],
reservoir_weight[68][85],
reservoir_weight[68][86],
reservoir_weight[68][87],
reservoir_weight[68][88],
reservoir_weight[68][89],
reservoir_weight[68][90],
reservoir_weight[68][91],
reservoir_weight[68][92],
reservoir_weight[68][93],
reservoir_weight[68][94],
reservoir_weight[68][95],
reservoir_weight[68][96],
reservoir_weight[68][97],
reservoir_weight[68][98],
reservoir_weight[68][99],
reservoir_weight[68][100],
reservoir_weight[68][101],
reservoir_weight[68][102],
reservoir_weight[68][103],
reservoir_weight[68][104],
reservoir_weight[68][105],
reservoir_weight[68][106],
reservoir_weight[68][107],
reservoir_weight[68][108],
reservoir_weight[68][109],
reservoir_weight[68][110],
reservoir_weight[68][111],
reservoir_weight[68][112],
reservoir_weight[68][113],
reservoir_weight[68][114],
reservoir_weight[68][115],
reservoir_weight[68][116],
reservoir_weight[68][117],
reservoir_weight[68][118],
reservoir_weight[68][119],
reservoir_weight[68][120],
reservoir_weight[68][121],
reservoir_weight[68][122],
reservoir_weight[68][123],
reservoir_weight[68][124],
reservoir_weight[68][125],
reservoir_weight[68][126],
reservoir_weight[68][127],
reservoir_weight[68][128],
reservoir_weight[68][129],
reservoir_weight[68][130],
reservoir_weight[68][131],
reservoir_weight[68][132],
reservoir_weight[68][133],
reservoir_weight[68][134],
reservoir_weight[68][135],
reservoir_weight[68][136],
reservoir_weight[68][137],
reservoir_weight[68][138],
reservoir_weight[68][139],
reservoir_weight[68][140],
reservoir_weight[68][141],
reservoir_weight[68][142],
reservoir_weight[68][143],
reservoir_weight[68][144],
reservoir_weight[68][145],
reservoir_weight[68][146],
reservoir_weight[68][147],
reservoir_weight[68][148],
reservoir_weight[68][149],
reservoir_weight[68][150],
reservoir_weight[68][151],
reservoir_weight[68][152],
reservoir_weight[68][153],
reservoir_weight[68][154],
reservoir_weight[68][155],
reservoir_weight[68][156],
reservoir_weight[68][157],
reservoir_weight[68][158],
reservoir_weight[68][159],
reservoir_weight[68][160],
reservoir_weight[68][161],
reservoir_weight[68][162],
reservoir_weight[68][163],
reservoir_weight[68][164],
reservoir_weight[68][165],
reservoir_weight[68][166],
reservoir_weight[68][167],
reservoir_weight[68][168],
reservoir_weight[68][169],
reservoir_weight[68][170],
reservoir_weight[68][171],
reservoir_weight[68][172],
reservoir_weight[68][173],
reservoir_weight[68][174],
reservoir_weight[68][175],
reservoir_weight[68][176],
reservoir_weight[68][177],
reservoir_weight[68][178],
reservoir_weight[68][179],
reservoir_weight[68][180],
reservoir_weight[68][181],
reservoir_weight[68][182],
reservoir_weight[68][183],
reservoir_weight[68][184],
reservoir_weight[68][185],
reservoir_weight[68][186],
reservoir_weight[68][187],
reservoir_weight[68][188],
reservoir_weight[68][189],
reservoir_weight[68][190],
reservoir_weight[68][191],
reservoir_weight[68][192],
reservoir_weight[68][193],
reservoir_weight[68][194],
reservoir_weight[68][195],
reservoir_weight[68][196],
reservoir_weight[68][197],
reservoir_weight[68][198],
reservoir_weight[68][199]
},
{reservoir_weight[69][0],
reservoir_weight[69][1],
reservoir_weight[69][2],
reservoir_weight[69][3],
reservoir_weight[69][4],
reservoir_weight[69][5],
reservoir_weight[69][6],
reservoir_weight[69][7],
reservoir_weight[69][8],
reservoir_weight[69][9],
reservoir_weight[69][10],
reservoir_weight[69][11],
reservoir_weight[69][12],
reservoir_weight[69][13],
reservoir_weight[69][14],
reservoir_weight[69][15],
reservoir_weight[69][16],
reservoir_weight[69][17],
reservoir_weight[69][18],
reservoir_weight[69][19],
reservoir_weight[69][20],
reservoir_weight[69][21],
reservoir_weight[69][22],
reservoir_weight[69][23],
reservoir_weight[69][24],
reservoir_weight[69][25],
reservoir_weight[69][26],
reservoir_weight[69][27],
reservoir_weight[69][28],
reservoir_weight[69][29],
reservoir_weight[69][30],
reservoir_weight[69][31],
reservoir_weight[69][32],
reservoir_weight[69][33],
reservoir_weight[69][34],
reservoir_weight[69][35],
reservoir_weight[69][36],
reservoir_weight[69][37],
reservoir_weight[69][38],
reservoir_weight[69][39],
reservoir_weight[69][40],
reservoir_weight[69][41],
reservoir_weight[69][42],
reservoir_weight[69][43],
reservoir_weight[69][44],
reservoir_weight[69][45],
reservoir_weight[69][46],
reservoir_weight[69][47],
reservoir_weight[69][48],
reservoir_weight[69][49],
reservoir_weight[69][50],
reservoir_weight[69][51],
reservoir_weight[69][52],
reservoir_weight[69][53],
reservoir_weight[69][54],
reservoir_weight[69][55],
reservoir_weight[69][56],
reservoir_weight[69][57],
reservoir_weight[69][58],
reservoir_weight[69][59],
reservoir_weight[69][60],
reservoir_weight[69][61],
reservoir_weight[69][62],
reservoir_weight[69][63],
reservoir_weight[69][64],
reservoir_weight[69][65],
reservoir_weight[69][66],
reservoir_weight[69][67],
reservoir_weight[69][68],
reservoir_weight[69][69],
reservoir_weight[69][70],
reservoir_weight[69][71],
reservoir_weight[69][72],
reservoir_weight[69][73],
reservoir_weight[69][74],
reservoir_weight[69][75],
reservoir_weight[69][76],
reservoir_weight[69][77],
reservoir_weight[69][78],
reservoir_weight[69][79],
reservoir_weight[69][80],
reservoir_weight[69][81],
reservoir_weight[69][82],
reservoir_weight[69][83],
reservoir_weight[69][84],
reservoir_weight[69][85],
reservoir_weight[69][86],
reservoir_weight[69][87],
reservoir_weight[69][88],
reservoir_weight[69][89],
reservoir_weight[69][90],
reservoir_weight[69][91],
reservoir_weight[69][92],
reservoir_weight[69][93],
reservoir_weight[69][94],
reservoir_weight[69][95],
reservoir_weight[69][96],
reservoir_weight[69][97],
reservoir_weight[69][98],
reservoir_weight[69][99],
reservoir_weight[69][100],
reservoir_weight[69][101],
reservoir_weight[69][102],
reservoir_weight[69][103],
reservoir_weight[69][104],
reservoir_weight[69][105],
reservoir_weight[69][106],
reservoir_weight[69][107],
reservoir_weight[69][108],
reservoir_weight[69][109],
reservoir_weight[69][110],
reservoir_weight[69][111],
reservoir_weight[69][112],
reservoir_weight[69][113],
reservoir_weight[69][114],
reservoir_weight[69][115],
reservoir_weight[69][116],
reservoir_weight[69][117],
reservoir_weight[69][118],
reservoir_weight[69][119],
reservoir_weight[69][120],
reservoir_weight[69][121],
reservoir_weight[69][122],
reservoir_weight[69][123],
reservoir_weight[69][124],
reservoir_weight[69][125],
reservoir_weight[69][126],
reservoir_weight[69][127],
reservoir_weight[69][128],
reservoir_weight[69][129],
reservoir_weight[69][130],
reservoir_weight[69][131],
reservoir_weight[69][132],
reservoir_weight[69][133],
reservoir_weight[69][134],
reservoir_weight[69][135],
reservoir_weight[69][136],
reservoir_weight[69][137],
reservoir_weight[69][138],
reservoir_weight[69][139],
reservoir_weight[69][140],
reservoir_weight[69][141],
reservoir_weight[69][142],
reservoir_weight[69][143],
reservoir_weight[69][144],
reservoir_weight[69][145],
reservoir_weight[69][146],
reservoir_weight[69][147],
reservoir_weight[69][148],
reservoir_weight[69][149],
reservoir_weight[69][150],
reservoir_weight[69][151],
reservoir_weight[69][152],
reservoir_weight[69][153],
reservoir_weight[69][154],
reservoir_weight[69][155],
reservoir_weight[69][156],
reservoir_weight[69][157],
reservoir_weight[69][158],
reservoir_weight[69][159],
reservoir_weight[69][160],
reservoir_weight[69][161],
reservoir_weight[69][162],
reservoir_weight[69][163],
reservoir_weight[69][164],
reservoir_weight[69][165],
reservoir_weight[69][166],
reservoir_weight[69][167],
reservoir_weight[69][168],
reservoir_weight[69][169],
reservoir_weight[69][170],
reservoir_weight[69][171],
reservoir_weight[69][172],
reservoir_weight[69][173],
reservoir_weight[69][174],
reservoir_weight[69][175],
reservoir_weight[69][176],
reservoir_weight[69][177],
reservoir_weight[69][178],
reservoir_weight[69][179],
reservoir_weight[69][180],
reservoir_weight[69][181],
reservoir_weight[69][182],
reservoir_weight[69][183],
reservoir_weight[69][184],
reservoir_weight[69][185],
reservoir_weight[69][186],
reservoir_weight[69][187],
reservoir_weight[69][188],
reservoir_weight[69][189],
reservoir_weight[69][190],
reservoir_weight[69][191],
reservoir_weight[69][192],
reservoir_weight[69][193],
reservoir_weight[69][194],
reservoir_weight[69][195],
reservoir_weight[69][196],
reservoir_weight[69][197],
reservoir_weight[69][198],
reservoir_weight[69][199]
},
{reservoir_weight[70][0],
reservoir_weight[70][1],
reservoir_weight[70][2],
reservoir_weight[70][3],
reservoir_weight[70][4],
reservoir_weight[70][5],
reservoir_weight[70][6],
reservoir_weight[70][7],
reservoir_weight[70][8],
reservoir_weight[70][9],
reservoir_weight[70][10],
reservoir_weight[70][11],
reservoir_weight[70][12],
reservoir_weight[70][13],
reservoir_weight[70][14],
reservoir_weight[70][15],
reservoir_weight[70][16],
reservoir_weight[70][17],
reservoir_weight[70][18],
reservoir_weight[70][19],
reservoir_weight[70][20],
reservoir_weight[70][21],
reservoir_weight[70][22],
reservoir_weight[70][23],
reservoir_weight[70][24],
reservoir_weight[70][25],
reservoir_weight[70][26],
reservoir_weight[70][27],
reservoir_weight[70][28],
reservoir_weight[70][29],
reservoir_weight[70][30],
reservoir_weight[70][31],
reservoir_weight[70][32],
reservoir_weight[70][33],
reservoir_weight[70][34],
reservoir_weight[70][35],
reservoir_weight[70][36],
reservoir_weight[70][37],
reservoir_weight[70][38],
reservoir_weight[70][39],
reservoir_weight[70][40],
reservoir_weight[70][41],
reservoir_weight[70][42],
reservoir_weight[70][43],
reservoir_weight[70][44],
reservoir_weight[70][45],
reservoir_weight[70][46],
reservoir_weight[70][47],
reservoir_weight[70][48],
reservoir_weight[70][49],
reservoir_weight[70][50],
reservoir_weight[70][51],
reservoir_weight[70][52],
reservoir_weight[70][53],
reservoir_weight[70][54],
reservoir_weight[70][55],
reservoir_weight[70][56],
reservoir_weight[70][57],
reservoir_weight[70][58],
reservoir_weight[70][59],
reservoir_weight[70][60],
reservoir_weight[70][61],
reservoir_weight[70][62],
reservoir_weight[70][63],
reservoir_weight[70][64],
reservoir_weight[70][65],
reservoir_weight[70][66],
reservoir_weight[70][67],
reservoir_weight[70][68],
reservoir_weight[70][69],
reservoir_weight[70][70],
reservoir_weight[70][71],
reservoir_weight[70][72],
reservoir_weight[70][73],
reservoir_weight[70][74],
reservoir_weight[70][75],
reservoir_weight[70][76],
reservoir_weight[70][77],
reservoir_weight[70][78],
reservoir_weight[70][79],
reservoir_weight[70][80],
reservoir_weight[70][81],
reservoir_weight[70][82],
reservoir_weight[70][83],
reservoir_weight[70][84],
reservoir_weight[70][85],
reservoir_weight[70][86],
reservoir_weight[70][87],
reservoir_weight[70][88],
reservoir_weight[70][89],
reservoir_weight[70][90],
reservoir_weight[70][91],
reservoir_weight[70][92],
reservoir_weight[70][93],
reservoir_weight[70][94],
reservoir_weight[70][95],
reservoir_weight[70][96],
reservoir_weight[70][97],
reservoir_weight[70][98],
reservoir_weight[70][99],
reservoir_weight[70][100],
reservoir_weight[70][101],
reservoir_weight[70][102],
reservoir_weight[70][103],
reservoir_weight[70][104],
reservoir_weight[70][105],
reservoir_weight[70][106],
reservoir_weight[70][107],
reservoir_weight[70][108],
reservoir_weight[70][109],
reservoir_weight[70][110],
reservoir_weight[70][111],
reservoir_weight[70][112],
reservoir_weight[70][113],
reservoir_weight[70][114],
reservoir_weight[70][115],
reservoir_weight[70][116],
reservoir_weight[70][117],
reservoir_weight[70][118],
reservoir_weight[70][119],
reservoir_weight[70][120],
reservoir_weight[70][121],
reservoir_weight[70][122],
reservoir_weight[70][123],
reservoir_weight[70][124],
reservoir_weight[70][125],
reservoir_weight[70][126],
reservoir_weight[70][127],
reservoir_weight[70][128],
reservoir_weight[70][129],
reservoir_weight[70][130],
reservoir_weight[70][131],
reservoir_weight[70][132],
reservoir_weight[70][133],
reservoir_weight[70][134],
reservoir_weight[70][135],
reservoir_weight[70][136],
reservoir_weight[70][137],
reservoir_weight[70][138],
reservoir_weight[70][139],
reservoir_weight[70][140],
reservoir_weight[70][141],
reservoir_weight[70][142],
reservoir_weight[70][143],
reservoir_weight[70][144],
reservoir_weight[70][145],
reservoir_weight[70][146],
reservoir_weight[70][147],
reservoir_weight[70][148],
reservoir_weight[70][149],
reservoir_weight[70][150],
reservoir_weight[70][151],
reservoir_weight[70][152],
reservoir_weight[70][153],
reservoir_weight[70][154],
reservoir_weight[70][155],
reservoir_weight[70][156],
reservoir_weight[70][157],
reservoir_weight[70][158],
reservoir_weight[70][159],
reservoir_weight[70][160],
reservoir_weight[70][161],
reservoir_weight[70][162],
reservoir_weight[70][163],
reservoir_weight[70][164],
reservoir_weight[70][165],
reservoir_weight[70][166],
reservoir_weight[70][167],
reservoir_weight[70][168],
reservoir_weight[70][169],
reservoir_weight[70][170],
reservoir_weight[70][171],
reservoir_weight[70][172],
reservoir_weight[70][173],
reservoir_weight[70][174],
reservoir_weight[70][175],
reservoir_weight[70][176],
reservoir_weight[70][177],
reservoir_weight[70][178],
reservoir_weight[70][179],
reservoir_weight[70][180],
reservoir_weight[70][181],
reservoir_weight[70][182],
reservoir_weight[70][183],
reservoir_weight[70][184],
reservoir_weight[70][185],
reservoir_weight[70][186],
reservoir_weight[70][187],
reservoir_weight[70][188],
reservoir_weight[70][189],
reservoir_weight[70][190],
reservoir_weight[70][191],
reservoir_weight[70][192],
reservoir_weight[70][193],
reservoir_weight[70][194],
reservoir_weight[70][195],
reservoir_weight[70][196],
reservoir_weight[70][197],
reservoir_weight[70][198],
reservoir_weight[70][199]
},
{reservoir_weight[71][0],
reservoir_weight[71][1],
reservoir_weight[71][2],
reservoir_weight[71][3],
reservoir_weight[71][4],
reservoir_weight[71][5],
reservoir_weight[71][6],
reservoir_weight[71][7],
reservoir_weight[71][8],
reservoir_weight[71][9],
reservoir_weight[71][10],
reservoir_weight[71][11],
reservoir_weight[71][12],
reservoir_weight[71][13],
reservoir_weight[71][14],
reservoir_weight[71][15],
reservoir_weight[71][16],
reservoir_weight[71][17],
reservoir_weight[71][18],
reservoir_weight[71][19],
reservoir_weight[71][20],
reservoir_weight[71][21],
reservoir_weight[71][22],
reservoir_weight[71][23],
reservoir_weight[71][24],
reservoir_weight[71][25],
reservoir_weight[71][26],
reservoir_weight[71][27],
reservoir_weight[71][28],
reservoir_weight[71][29],
reservoir_weight[71][30],
reservoir_weight[71][31],
reservoir_weight[71][32],
reservoir_weight[71][33],
reservoir_weight[71][34],
reservoir_weight[71][35],
reservoir_weight[71][36],
reservoir_weight[71][37],
reservoir_weight[71][38],
reservoir_weight[71][39],
reservoir_weight[71][40],
reservoir_weight[71][41],
reservoir_weight[71][42],
reservoir_weight[71][43],
reservoir_weight[71][44],
reservoir_weight[71][45],
reservoir_weight[71][46],
reservoir_weight[71][47],
reservoir_weight[71][48],
reservoir_weight[71][49],
reservoir_weight[71][50],
reservoir_weight[71][51],
reservoir_weight[71][52],
reservoir_weight[71][53],
reservoir_weight[71][54],
reservoir_weight[71][55],
reservoir_weight[71][56],
reservoir_weight[71][57],
reservoir_weight[71][58],
reservoir_weight[71][59],
reservoir_weight[71][60],
reservoir_weight[71][61],
reservoir_weight[71][62],
reservoir_weight[71][63],
reservoir_weight[71][64],
reservoir_weight[71][65],
reservoir_weight[71][66],
reservoir_weight[71][67],
reservoir_weight[71][68],
reservoir_weight[71][69],
reservoir_weight[71][70],
reservoir_weight[71][71],
reservoir_weight[71][72],
reservoir_weight[71][73],
reservoir_weight[71][74],
reservoir_weight[71][75],
reservoir_weight[71][76],
reservoir_weight[71][77],
reservoir_weight[71][78],
reservoir_weight[71][79],
reservoir_weight[71][80],
reservoir_weight[71][81],
reservoir_weight[71][82],
reservoir_weight[71][83],
reservoir_weight[71][84],
reservoir_weight[71][85],
reservoir_weight[71][86],
reservoir_weight[71][87],
reservoir_weight[71][88],
reservoir_weight[71][89],
reservoir_weight[71][90],
reservoir_weight[71][91],
reservoir_weight[71][92],
reservoir_weight[71][93],
reservoir_weight[71][94],
reservoir_weight[71][95],
reservoir_weight[71][96],
reservoir_weight[71][97],
reservoir_weight[71][98],
reservoir_weight[71][99],
reservoir_weight[71][100],
reservoir_weight[71][101],
reservoir_weight[71][102],
reservoir_weight[71][103],
reservoir_weight[71][104],
reservoir_weight[71][105],
reservoir_weight[71][106],
reservoir_weight[71][107],
reservoir_weight[71][108],
reservoir_weight[71][109],
reservoir_weight[71][110],
reservoir_weight[71][111],
reservoir_weight[71][112],
reservoir_weight[71][113],
reservoir_weight[71][114],
reservoir_weight[71][115],
reservoir_weight[71][116],
reservoir_weight[71][117],
reservoir_weight[71][118],
reservoir_weight[71][119],
reservoir_weight[71][120],
reservoir_weight[71][121],
reservoir_weight[71][122],
reservoir_weight[71][123],
reservoir_weight[71][124],
reservoir_weight[71][125],
reservoir_weight[71][126],
reservoir_weight[71][127],
reservoir_weight[71][128],
reservoir_weight[71][129],
reservoir_weight[71][130],
reservoir_weight[71][131],
reservoir_weight[71][132],
reservoir_weight[71][133],
reservoir_weight[71][134],
reservoir_weight[71][135],
reservoir_weight[71][136],
reservoir_weight[71][137],
reservoir_weight[71][138],
reservoir_weight[71][139],
reservoir_weight[71][140],
reservoir_weight[71][141],
reservoir_weight[71][142],
reservoir_weight[71][143],
reservoir_weight[71][144],
reservoir_weight[71][145],
reservoir_weight[71][146],
reservoir_weight[71][147],
reservoir_weight[71][148],
reservoir_weight[71][149],
reservoir_weight[71][150],
reservoir_weight[71][151],
reservoir_weight[71][152],
reservoir_weight[71][153],
reservoir_weight[71][154],
reservoir_weight[71][155],
reservoir_weight[71][156],
reservoir_weight[71][157],
reservoir_weight[71][158],
reservoir_weight[71][159],
reservoir_weight[71][160],
reservoir_weight[71][161],
reservoir_weight[71][162],
reservoir_weight[71][163],
reservoir_weight[71][164],
reservoir_weight[71][165],
reservoir_weight[71][166],
reservoir_weight[71][167],
reservoir_weight[71][168],
reservoir_weight[71][169],
reservoir_weight[71][170],
reservoir_weight[71][171],
reservoir_weight[71][172],
reservoir_weight[71][173],
reservoir_weight[71][174],
reservoir_weight[71][175],
reservoir_weight[71][176],
reservoir_weight[71][177],
reservoir_weight[71][178],
reservoir_weight[71][179],
reservoir_weight[71][180],
reservoir_weight[71][181],
reservoir_weight[71][182],
reservoir_weight[71][183],
reservoir_weight[71][184],
reservoir_weight[71][185],
reservoir_weight[71][186],
reservoir_weight[71][187],
reservoir_weight[71][188],
reservoir_weight[71][189],
reservoir_weight[71][190],
reservoir_weight[71][191],
reservoir_weight[71][192],
reservoir_weight[71][193],
reservoir_weight[71][194],
reservoir_weight[71][195],
reservoir_weight[71][196],
reservoir_weight[71][197],
reservoir_weight[71][198],
reservoir_weight[71][199]
},
{reservoir_weight[72][0],
reservoir_weight[72][1],
reservoir_weight[72][2],
reservoir_weight[72][3],
reservoir_weight[72][4],
reservoir_weight[72][5],
reservoir_weight[72][6],
reservoir_weight[72][7],
reservoir_weight[72][8],
reservoir_weight[72][9],
reservoir_weight[72][10],
reservoir_weight[72][11],
reservoir_weight[72][12],
reservoir_weight[72][13],
reservoir_weight[72][14],
reservoir_weight[72][15],
reservoir_weight[72][16],
reservoir_weight[72][17],
reservoir_weight[72][18],
reservoir_weight[72][19],
reservoir_weight[72][20],
reservoir_weight[72][21],
reservoir_weight[72][22],
reservoir_weight[72][23],
reservoir_weight[72][24],
reservoir_weight[72][25],
reservoir_weight[72][26],
reservoir_weight[72][27],
reservoir_weight[72][28],
reservoir_weight[72][29],
reservoir_weight[72][30],
reservoir_weight[72][31],
reservoir_weight[72][32],
reservoir_weight[72][33],
reservoir_weight[72][34],
reservoir_weight[72][35],
reservoir_weight[72][36],
reservoir_weight[72][37],
reservoir_weight[72][38],
reservoir_weight[72][39],
reservoir_weight[72][40],
reservoir_weight[72][41],
reservoir_weight[72][42],
reservoir_weight[72][43],
reservoir_weight[72][44],
reservoir_weight[72][45],
reservoir_weight[72][46],
reservoir_weight[72][47],
reservoir_weight[72][48],
reservoir_weight[72][49],
reservoir_weight[72][50],
reservoir_weight[72][51],
reservoir_weight[72][52],
reservoir_weight[72][53],
reservoir_weight[72][54],
reservoir_weight[72][55],
reservoir_weight[72][56],
reservoir_weight[72][57],
reservoir_weight[72][58],
reservoir_weight[72][59],
reservoir_weight[72][60],
reservoir_weight[72][61],
reservoir_weight[72][62],
reservoir_weight[72][63],
reservoir_weight[72][64],
reservoir_weight[72][65],
reservoir_weight[72][66],
reservoir_weight[72][67],
reservoir_weight[72][68],
reservoir_weight[72][69],
reservoir_weight[72][70],
reservoir_weight[72][71],
reservoir_weight[72][72],
reservoir_weight[72][73],
reservoir_weight[72][74],
reservoir_weight[72][75],
reservoir_weight[72][76],
reservoir_weight[72][77],
reservoir_weight[72][78],
reservoir_weight[72][79],
reservoir_weight[72][80],
reservoir_weight[72][81],
reservoir_weight[72][82],
reservoir_weight[72][83],
reservoir_weight[72][84],
reservoir_weight[72][85],
reservoir_weight[72][86],
reservoir_weight[72][87],
reservoir_weight[72][88],
reservoir_weight[72][89],
reservoir_weight[72][90],
reservoir_weight[72][91],
reservoir_weight[72][92],
reservoir_weight[72][93],
reservoir_weight[72][94],
reservoir_weight[72][95],
reservoir_weight[72][96],
reservoir_weight[72][97],
reservoir_weight[72][98],
reservoir_weight[72][99],
reservoir_weight[72][100],
reservoir_weight[72][101],
reservoir_weight[72][102],
reservoir_weight[72][103],
reservoir_weight[72][104],
reservoir_weight[72][105],
reservoir_weight[72][106],
reservoir_weight[72][107],
reservoir_weight[72][108],
reservoir_weight[72][109],
reservoir_weight[72][110],
reservoir_weight[72][111],
reservoir_weight[72][112],
reservoir_weight[72][113],
reservoir_weight[72][114],
reservoir_weight[72][115],
reservoir_weight[72][116],
reservoir_weight[72][117],
reservoir_weight[72][118],
reservoir_weight[72][119],
reservoir_weight[72][120],
reservoir_weight[72][121],
reservoir_weight[72][122],
reservoir_weight[72][123],
reservoir_weight[72][124],
reservoir_weight[72][125],
reservoir_weight[72][126],
reservoir_weight[72][127],
reservoir_weight[72][128],
reservoir_weight[72][129],
reservoir_weight[72][130],
reservoir_weight[72][131],
reservoir_weight[72][132],
reservoir_weight[72][133],
reservoir_weight[72][134],
reservoir_weight[72][135],
reservoir_weight[72][136],
reservoir_weight[72][137],
reservoir_weight[72][138],
reservoir_weight[72][139],
reservoir_weight[72][140],
reservoir_weight[72][141],
reservoir_weight[72][142],
reservoir_weight[72][143],
reservoir_weight[72][144],
reservoir_weight[72][145],
reservoir_weight[72][146],
reservoir_weight[72][147],
reservoir_weight[72][148],
reservoir_weight[72][149],
reservoir_weight[72][150],
reservoir_weight[72][151],
reservoir_weight[72][152],
reservoir_weight[72][153],
reservoir_weight[72][154],
reservoir_weight[72][155],
reservoir_weight[72][156],
reservoir_weight[72][157],
reservoir_weight[72][158],
reservoir_weight[72][159],
reservoir_weight[72][160],
reservoir_weight[72][161],
reservoir_weight[72][162],
reservoir_weight[72][163],
reservoir_weight[72][164],
reservoir_weight[72][165],
reservoir_weight[72][166],
reservoir_weight[72][167],
reservoir_weight[72][168],
reservoir_weight[72][169],
reservoir_weight[72][170],
reservoir_weight[72][171],
reservoir_weight[72][172],
reservoir_weight[72][173],
reservoir_weight[72][174],
reservoir_weight[72][175],
reservoir_weight[72][176],
reservoir_weight[72][177],
reservoir_weight[72][178],
reservoir_weight[72][179],
reservoir_weight[72][180],
reservoir_weight[72][181],
reservoir_weight[72][182],
reservoir_weight[72][183],
reservoir_weight[72][184],
reservoir_weight[72][185],
reservoir_weight[72][186],
reservoir_weight[72][187],
reservoir_weight[72][188],
reservoir_weight[72][189],
reservoir_weight[72][190],
reservoir_weight[72][191],
reservoir_weight[72][192],
reservoir_weight[72][193],
reservoir_weight[72][194],
reservoir_weight[72][195],
reservoir_weight[72][196],
reservoir_weight[72][197],
reservoir_weight[72][198],
reservoir_weight[72][199]
},
{reservoir_weight[73][0],
reservoir_weight[73][1],
reservoir_weight[73][2],
reservoir_weight[73][3],
reservoir_weight[73][4],
reservoir_weight[73][5],
reservoir_weight[73][6],
reservoir_weight[73][7],
reservoir_weight[73][8],
reservoir_weight[73][9],
reservoir_weight[73][10],
reservoir_weight[73][11],
reservoir_weight[73][12],
reservoir_weight[73][13],
reservoir_weight[73][14],
reservoir_weight[73][15],
reservoir_weight[73][16],
reservoir_weight[73][17],
reservoir_weight[73][18],
reservoir_weight[73][19],
reservoir_weight[73][20],
reservoir_weight[73][21],
reservoir_weight[73][22],
reservoir_weight[73][23],
reservoir_weight[73][24],
reservoir_weight[73][25],
reservoir_weight[73][26],
reservoir_weight[73][27],
reservoir_weight[73][28],
reservoir_weight[73][29],
reservoir_weight[73][30],
reservoir_weight[73][31],
reservoir_weight[73][32],
reservoir_weight[73][33],
reservoir_weight[73][34],
reservoir_weight[73][35],
reservoir_weight[73][36],
reservoir_weight[73][37],
reservoir_weight[73][38],
reservoir_weight[73][39],
reservoir_weight[73][40],
reservoir_weight[73][41],
reservoir_weight[73][42],
reservoir_weight[73][43],
reservoir_weight[73][44],
reservoir_weight[73][45],
reservoir_weight[73][46],
reservoir_weight[73][47],
reservoir_weight[73][48],
reservoir_weight[73][49],
reservoir_weight[73][50],
reservoir_weight[73][51],
reservoir_weight[73][52],
reservoir_weight[73][53],
reservoir_weight[73][54],
reservoir_weight[73][55],
reservoir_weight[73][56],
reservoir_weight[73][57],
reservoir_weight[73][58],
reservoir_weight[73][59],
reservoir_weight[73][60],
reservoir_weight[73][61],
reservoir_weight[73][62],
reservoir_weight[73][63],
reservoir_weight[73][64],
reservoir_weight[73][65],
reservoir_weight[73][66],
reservoir_weight[73][67],
reservoir_weight[73][68],
reservoir_weight[73][69],
reservoir_weight[73][70],
reservoir_weight[73][71],
reservoir_weight[73][72],
reservoir_weight[73][73],
reservoir_weight[73][74],
reservoir_weight[73][75],
reservoir_weight[73][76],
reservoir_weight[73][77],
reservoir_weight[73][78],
reservoir_weight[73][79],
reservoir_weight[73][80],
reservoir_weight[73][81],
reservoir_weight[73][82],
reservoir_weight[73][83],
reservoir_weight[73][84],
reservoir_weight[73][85],
reservoir_weight[73][86],
reservoir_weight[73][87],
reservoir_weight[73][88],
reservoir_weight[73][89],
reservoir_weight[73][90],
reservoir_weight[73][91],
reservoir_weight[73][92],
reservoir_weight[73][93],
reservoir_weight[73][94],
reservoir_weight[73][95],
reservoir_weight[73][96],
reservoir_weight[73][97],
reservoir_weight[73][98],
reservoir_weight[73][99],
reservoir_weight[73][100],
reservoir_weight[73][101],
reservoir_weight[73][102],
reservoir_weight[73][103],
reservoir_weight[73][104],
reservoir_weight[73][105],
reservoir_weight[73][106],
reservoir_weight[73][107],
reservoir_weight[73][108],
reservoir_weight[73][109],
reservoir_weight[73][110],
reservoir_weight[73][111],
reservoir_weight[73][112],
reservoir_weight[73][113],
reservoir_weight[73][114],
reservoir_weight[73][115],
reservoir_weight[73][116],
reservoir_weight[73][117],
reservoir_weight[73][118],
reservoir_weight[73][119],
reservoir_weight[73][120],
reservoir_weight[73][121],
reservoir_weight[73][122],
reservoir_weight[73][123],
reservoir_weight[73][124],
reservoir_weight[73][125],
reservoir_weight[73][126],
reservoir_weight[73][127],
reservoir_weight[73][128],
reservoir_weight[73][129],
reservoir_weight[73][130],
reservoir_weight[73][131],
reservoir_weight[73][132],
reservoir_weight[73][133],
reservoir_weight[73][134],
reservoir_weight[73][135],
reservoir_weight[73][136],
reservoir_weight[73][137],
reservoir_weight[73][138],
reservoir_weight[73][139],
reservoir_weight[73][140],
reservoir_weight[73][141],
reservoir_weight[73][142],
reservoir_weight[73][143],
reservoir_weight[73][144],
reservoir_weight[73][145],
reservoir_weight[73][146],
reservoir_weight[73][147],
reservoir_weight[73][148],
reservoir_weight[73][149],
reservoir_weight[73][150],
reservoir_weight[73][151],
reservoir_weight[73][152],
reservoir_weight[73][153],
reservoir_weight[73][154],
reservoir_weight[73][155],
reservoir_weight[73][156],
reservoir_weight[73][157],
reservoir_weight[73][158],
reservoir_weight[73][159],
reservoir_weight[73][160],
reservoir_weight[73][161],
reservoir_weight[73][162],
reservoir_weight[73][163],
reservoir_weight[73][164],
reservoir_weight[73][165],
reservoir_weight[73][166],
reservoir_weight[73][167],
reservoir_weight[73][168],
reservoir_weight[73][169],
reservoir_weight[73][170],
reservoir_weight[73][171],
reservoir_weight[73][172],
reservoir_weight[73][173],
reservoir_weight[73][174],
reservoir_weight[73][175],
reservoir_weight[73][176],
reservoir_weight[73][177],
reservoir_weight[73][178],
reservoir_weight[73][179],
reservoir_weight[73][180],
reservoir_weight[73][181],
reservoir_weight[73][182],
reservoir_weight[73][183],
reservoir_weight[73][184],
reservoir_weight[73][185],
reservoir_weight[73][186],
reservoir_weight[73][187],
reservoir_weight[73][188],
reservoir_weight[73][189],
reservoir_weight[73][190],
reservoir_weight[73][191],
reservoir_weight[73][192],
reservoir_weight[73][193],
reservoir_weight[73][194],
reservoir_weight[73][195],
reservoir_weight[73][196],
reservoir_weight[73][197],
reservoir_weight[73][198],
reservoir_weight[73][199]
},
{reservoir_weight[74][0],
reservoir_weight[74][1],
reservoir_weight[74][2],
reservoir_weight[74][3],
reservoir_weight[74][4],
reservoir_weight[74][5],
reservoir_weight[74][6],
reservoir_weight[74][7],
reservoir_weight[74][8],
reservoir_weight[74][9],
reservoir_weight[74][10],
reservoir_weight[74][11],
reservoir_weight[74][12],
reservoir_weight[74][13],
reservoir_weight[74][14],
reservoir_weight[74][15],
reservoir_weight[74][16],
reservoir_weight[74][17],
reservoir_weight[74][18],
reservoir_weight[74][19],
reservoir_weight[74][20],
reservoir_weight[74][21],
reservoir_weight[74][22],
reservoir_weight[74][23],
reservoir_weight[74][24],
reservoir_weight[74][25],
reservoir_weight[74][26],
reservoir_weight[74][27],
reservoir_weight[74][28],
reservoir_weight[74][29],
reservoir_weight[74][30],
reservoir_weight[74][31],
reservoir_weight[74][32],
reservoir_weight[74][33],
reservoir_weight[74][34],
reservoir_weight[74][35],
reservoir_weight[74][36],
reservoir_weight[74][37],
reservoir_weight[74][38],
reservoir_weight[74][39],
reservoir_weight[74][40],
reservoir_weight[74][41],
reservoir_weight[74][42],
reservoir_weight[74][43],
reservoir_weight[74][44],
reservoir_weight[74][45],
reservoir_weight[74][46],
reservoir_weight[74][47],
reservoir_weight[74][48],
reservoir_weight[74][49],
reservoir_weight[74][50],
reservoir_weight[74][51],
reservoir_weight[74][52],
reservoir_weight[74][53],
reservoir_weight[74][54],
reservoir_weight[74][55],
reservoir_weight[74][56],
reservoir_weight[74][57],
reservoir_weight[74][58],
reservoir_weight[74][59],
reservoir_weight[74][60],
reservoir_weight[74][61],
reservoir_weight[74][62],
reservoir_weight[74][63],
reservoir_weight[74][64],
reservoir_weight[74][65],
reservoir_weight[74][66],
reservoir_weight[74][67],
reservoir_weight[74][68],
reservoir_weight[74][69],
reservoir_weight[74][70],
reservoir_weight[74][71],
reservoir_weight[74][72],
reservoir_weight[74][73],
reservoir_weight[74][74],
reservoir_weight[74][75],
reservoir_weight[74][76],
reservoir_weight[74][77],
reservoir_weight[74][78],
reservoir_weight[74][79],
reservoir_weight[74][80],
reservoir_weight[74][81],
reservoir_weight[74][82],
reservoir_weight[74][83],
reservoir_weight[74][84],
reservoir_weight[74][85],
reservoir_weight[74][86],
reservoir_weight[74][87],
reservoir_weight[74][88],
reservoir_weight[74][89],
reservoir_weight[74][90],
reservoir_weight[74][91],
reservoir_weight[74][92],
reservoir_weight[74][93],
reservoir_weight[74][94],
reservoir_weight[74][95],
reservoir_weight[74][96],
reservoir_weight[74][97],
reservoir_weight[74][98],
reservoir_weight[74][99],
reservoir_weight[74][100],
reservoir_weight[74][101],
reservoir_weight[74][102],
reservoir_weight[74][103],
reservoir_weight[74][104],
reservoir_weight[74][105],
reservoir_weight[74][106],
reservoir_weight[74][107],
reservoir_weight[74][108],
reservoir_weight[74][109],
reservoir_weight[74][110],
reservoir_weight[74][111],
reservoir_weight[74][112],
reservoir_weight[74][113],
reservoir_weight[74][114],
reservoir_weight[74][115],
reservoir_weight[74][116],
reservoir_weight[74][117],
reservoir_weight[74][118],
reservoir_weight[74][119],
reservoir_weight[74][120],
reservoir_weight[74][121],
reservoir_weight[74][122],
reservoir_weight[74][123],
reservoir_weight[74][124],
reservoir_weight[74][125],
reservoir_weight[74][126],
reservoir_weight[74][127],
reservoir_weight[74][128],
reservoir_weight[74][129],
reservoir_weight[74][130],
reservoir_weight[74][131],
reservoir_weight[74][132],
reservoir_weight[74][133],
reservoir_weight[74][134],
reservoir_weight[74][135],
reservoir_weight[74][136],
reservoir_weight[74][137],
reservoir_weight[74][138],
reservoir_weight[74][139],
reservoir_weight[74][140],
reservoir_weight[74][141],
reservoir_weight[74][142],
reservoir_weight[74][143],
reservoir_weight[74][144],
reservoir_weight[74][145],
reservoir_weight[74][146],
reservoir_weight[74][147],
reservoir_weight[74][148],
reservoir_weight[74][149],
reservoir_weight[74][150],
reservoir_weight[74][151],
reservoir_weight[74][152],
reservoir_weight[74][153],
reservoir_weight[74][154],
reservoir_weight[74][155],
reservoir_weight[74][156],
reservoir_weight[74][157],
reservoir_weight[74][158],
reservoir_weight[74][159],
reservoir_weight[74][160],
reservoir_weight[74][161],
reservoir_weight[74][162],
reservoir_weight[74][163],
reservoir_weight[74][164],
reservoir_weight[74][165],
reservoir_weight[74][166],
reservoir_weight[74][167],
reservoir_weight[74][168],
reservoir_weight[74][169],
reservoir_weight[74][170],
reservoir_weight[74][171],
reservoir_weight[74][172],
reservoir_weight[74][173],
reservoir_weight[74][174],
reservoir_weight[74][175],
reservoir_weight[74][176],
reservoir_weight[74][177],
reservoir_weight[74][178],
reservoir_weight[74][179],
reservoir_weight[74][180],
reservoir_weight[74][181],
reservoir_weight[74][182],
reservoir_weight[74][183],
reservoir_weight[74][184],
reservoir_weight[74][185],
reservoir_weight[74][186],
reservoir_weight[74][187],
reservoir_weight[74][188],
reservoir_weight[74][189],
reservoir_weight[74][190],
reservoir_weight[74][191],
reservoir_weight[74][192],
reservoir_weight[74][193],
reservoir_weight[74][194],
reservoir_weight[74][195],
reservoir_weight[74][196],
reservoir_weight[74][197],
reservoir_weight[74][198],
reservoir_weight[74][199]
},
{reservoir_weight[75][0],
reservoir_weight[75][1],
reservoir_weight[75][2],
reservoir_weight[75][3],
reservoir_weight[75][4],
reservoir_weight[75][5],
reservoir_weight[75][6],
reservoir_weight[75][7],
reservoir_weight[75][8],
reservoir_weight[75][9],
reservoir_weight[75][10],
reservoir_weight[75][11],
reservoir_weight[75][12],
reservoir_weight[75][13],
reservoir_weight[75][14],
reservoir_weight[75][15],
reservoir_weight[75][16],
reservoir_weight[75][17],
reservoir_weight[75][18],
reservoir_weight[75][19],
reservoir_weight[75][20],
reservoir_weight[75][21],
reservoir_weight[75][22],
reservoir_weight[75][23],
reservoir_weight[75][24],
reservoir_weight[75][25],
reservoir_weight[75][26],
reservoir_weight[75][27],
reservoir_weight[75][28],
reservoir_weight[75][29],
reservoir_weight[75][30],
reservoir_weight[75][31],
reservoir_weight[75][32],
reservoir_weight[75][33],
reservoir_weight[75][34],
reservoir_weight[75][35],
reservoir_weight[75][36],
reservoir_weight[75][37],
reservoir_weight[75][38],
reservoir_weight[75][39],
reservoir_weight[75][40],
reservoir_weight[75][41],
reservoir_weight[75][42],
reservoir_weight[75][43],
reservoir_weight[75][44],
reservoir_weight[75][45],
reservoir_weight[75][46],
reservoir_weight[75][47],
reservoir_weight[75][48],
reservoir_weight[75][49],
reservoir_weight[75][50],
reservoir_weight[75][51],
reservoir_weight[75][52],
reservoir_weight[75][53],
reservoir_weight[75][54],
reservoir_weight[75][55],
reservoir_weight[75][56],
reservoir_weight[75][57],
reservoir_weight[75][58],
reservoir_weight[75][59],
reservoir_weight[75][60],
reservoir_weight[75][61],
reservoir_weight[75][62],
reservoir_weight[75][63],
reservoir_weight[75][64],
reservoir_weight[75][65],
reservoir_weight[75][66],
reservoir_weight[75][67],
reservoir_weight[75][68],
reservoir_weight[75][69],
reservoir_weight[75][70],
reservoir_weight[75][71],
reservoir_weight[75][72],
reservoir_weight[75][73],
reservoir_weight[75][74],
reservoir_weight[75][75],
reservoir_weight[75][76],
reservoir_weight[75][77],
reservoir_weight[75][78],
reservoir_weight[75][79],
reservoir_weight[75][80],
reservoir_weight[75][81],
reservoir_weight[75][82],
reservoir_weight[75][83],
reservoir_weight[75][84],
reservoir_weight[75][85],
reservoir_weight[75][86],
reservoir_weight[75][87],
reservoir_weight[75][88],
reservoir_weight[75][89],
reservoir_weight[75][90],
reservoir_weight[75][91],
reservoir_weight[75][92],
reservoir_weight[75][93],
reservoir_weight[75][94],
reservoir_weight[75][95],
reservoir_weight[75][96],
reservoir_weight[75][97],
reservoir_weight[75][98],
reservoir_weight[75][99],
reservoir_weight[75][100],
reservoir_weight[75][101],
reservoir_weight[75][102],
reservoir_weight[75][103],
reservoir_weight[75][104],
reservoir_weight[75][105],
reservoir_weight[75][106],
reservoir_weight[75][107],
reservoir_weight[75][108],
reservoir_weight[75][109],
reservoir_weight[75][110],
reservoir_weight[75][111],
reservoir_weight[75][112],
reservoir_weight[75][113],
reservoir_weight[75][114],
reservoir_weight[75][115],
reservoir_weight[75][116],
reservoir_weight[75][117],
reservoir_weight[75][118],
reservoir_weight[75][119],
reservoir_weight[75][120],
reservoir_weight[75][121],
reservoir_weight[75][122],
reservoir_weight[75][123],
reservoir_weight[75][124],
reservoir_weight[75][125],
reservoir_weight[75][126],
reservoir_weight[75][127],
reservoir_weight[75][128],
reservoir_weight[75][129],
reservoir_weight[75][130],
reservoir_weight[75][131],
reservoir_weight[75][132],
reservoir_weight[75][133],
reservoir_weight[75][134],
reservoir_weight[75][135],
reservoir_weight[75][136],
reservoir_weight[75][137],
reservoir_weight[75][138],
reservoir_weight[75][139],
reservoir_weight[75][140],
reservoir_weight[75][141],
reservoir_weight[75][142],
reservoir_weight[75][143],
reservoir_weight[75][144],
reservoir_weight[75][145],
reservoir_weight[75][146],
reservoir_weight[75][147],
reservoir_weight[75][148],
reservoir_weight[75][149],
reservoir_weight[75][150],
reservoir_weight[75][151],
reservoir_weight[75][152],
reservoir_weight[75][153],
reservoir_weight[75][154],
reservoir_weight[75][155],
reservoir_weight[75][156],
reservoir_weight[75][157],
reservoir_weight[75][158],
reservoir_weight[75][159],
reservoir_weight[75][160],
reservoir_weight[75][161],
reservoir_weight[75][162],
reservoir_weight[75][163],
reservoir_weight[75][164],
reservoir_weight[75][165],
reservoir_weight[75][166],
reservoir_weight[75][167],
reservoir_weight[75][168],
reservoir_weight[75][169],
reservoir_weight[75][170],
reservoir_weight[75][171],
reservoir_weight[75][172],
reservoir_weight[75][173],
reservoir_weight[75][174],
reservoir_weight[75][175],
reservoir_weight[75][176],
reservoir_weight[75][177],
reservoir_weight[75][178],
reservoir_weight[75][179],
reservoir_weight[75][180],
reservoir_weight[75][181],
reservoir_weight[75][182],
reservoir_weight[75][183],
reservoir_weight[75][184],
reservoir_weight[75][185],
reservoir_weight[75][186],
reservoir_weight[75][187],
reservoir_weight[75][188],
reservoir_weight[75][189],
reservoir_weight[75][190],
reservoir_weight[75][191],
reservoir_weight[75][192],
reservoir_weight[75][193],
reservoir_weight[75][194],
reservoir_weight[75][195],
reservoir_weight[75][196],
reservoir_weight[75][197],
reservoir_weight[75][198],
reservoir_weight[75][199]
},
{reservoir_weight[76][0],
reservoir_weight[76][1],
reservoir_weight[76][2],
reservoir_weight[76][3],
reservoir_weight[76][4],
reservoir_weight[76][5],
reservoir_weight[76][6],
reservoir_weight[76][7],
reservoir_weight[76][8],
reservoir_weight[76][9],
reservoir_weight[76][10],
reservoir_weight[76][11],
reservoir_weight[76][12],
reservoir_weight[76][13],
reservoir_weight[76][14],
reservoir_weight[76][15],
reservoir_weight[76][16],
reservoir_weight[76][17],
reservoir_weight[76][18],
reservoir_weight[76][19],
reservoir_weight[76][20],
reservoir_weight[76][21],
reservoir_weight[76][22],
reservoir_weight[76][23],
reservoir_weight[76][24],
reservoir_weight[76][25],
reservoir_weight[76][26],
reservoir_weight[76][27],
reservoir_weight[76][28],
reservoir_weight[76][29],
reservoir_weight[76][30],
reservoir_weight[76][31],
reservoir_weight[76][32],
reservoir_weight[76][33],
reservoir_weight[76][34],
reservoir_weight[76][35],
reservoir_weight[76][36],
reservoir_weight[76][37],
reservoir_weight[76][38],
reservoir_weight[76][39],
reservoir_weight[76][40],
reservoir_weight[76][41],
reservoir_weight[76][42],
reservoir_weight[76][43],
reservoir_weight[76][44],
reservoir_weight[76][45],
reservoir_weight[76][46],
reservoir_weight[76][47],
reservoir_weight[76][48],
reservoir_weight[76][49],
reservoir_weight[76][50],
reservoir_weight[76][51],
reservoir_weight[76][52],
reservoir_weight[76][53],
reservoir_weight[76][54],
reservoir_weight[76][55],
reservoir_weight[76][56],
reservoir_weight[76][57],
reservoir_weight[76][58],
reservoir_weight[76][59],
reservoir_weight[76][60],
reservoir_weight[76][61],
reservoir_weight[76][62],
reservoir_weight[76][63],
reservoir_weight[76][64],
reservoir_weight[76][65],
reservoir_weight[76][66],
reservoir_weight[76][67],
reservoir_weight[76][68],
reservoir_weight[76][69],
reservoir_weight[76][70],
reservoir_weight[76][71],
reservoir_weight[76][72],
reservoir_weight[76][73],
reservoir_weight[76][74],
reservoir_weight[76][75],
reservoir_weight[76][76],
reservoir_weight[76][77],
reservoir_weight[76][78],
reservoir_weight[76][79],
reservoir_weight[76][80],
reservoir_weight[76][81],
reservoir_weight[76][82],
reservoir_weight[76][83],
reservoir_weight[76][84],
reservoir_weight[76][85],
reservoir_weight[76][86],
reservoir_weight[76][87],
reservoir_weight[76][88],
reservoir_weight[76][89],
reservoir_weight[76][90],
reservoir_weight[76][91],
reservoir_weight[76][92],
reservoir_weight[76][93],
reservoir_weight[76][94],
reservoir_weight[76][95],
reservoir_weight[76][96],
reservoir_weight[76][97],
reservoir_weight[76][98],
reservoir_weight[76][99],
reservoir_weight[76][100],
reservoir_weight[76][101],
reservoir_weight[76][102],
reservoir_weight[76][103],
reservoir_weight[76][104],
reservoir_weight[76][105],
reservoir_weight[76][106],
reservoir_weight[76][107],
reservoir_weight[76][108],
reservoir_weight[76][109],
reservoir_weight[76][110],
reservoir_weight[76][111],
reservoir_weight[76][112],
reservoir_weight[76][113],
reservoir_weight[76][114],
reservoir_weight[76][115],
reservoir_weight[76][116],
reservoir_weight[76][117],
reservoir_weight[76][118],
reservoir_weight[76][119],
reservoir_weight[76][120],
reservoir_weight[76][121],
reservoir_weight[76][122],
reservoir_weight[76][123],
reservoir_weight[76][124],
reservoir_weight[76][125],
reservoir_weight[76][126],
reservoir_weight[76][127],
reservoir_weight[76][128],
reservoir_weight[76][129],
reservoir_weight[76][130],
reservoir_weight[76][131],
reservoir_weight[76][132],
reservoir_weight[76][133],
reservoir_weight[76][134],
reservoir_weight[76][135],
reservoir_weight[76][136],
reservoir_weight[76][137],
reservoir_weight[76][138],
reservoir_weight[76][139],
reservoir_weight[76][140],
reservoir_weight[76][141],
reservoir_weight[76][142],
reservoir_weight[76][143],
reservoir_weight[76][144],
reservoir_weight[76][145],
reservoir_weight[76][146],
reservoir_weight[76][147],
reservoir_weight[76][148],
reservoir_weight[76][149],
reservoir_weight[76][150],
reservoir_weight[76][151],
reservoir_weight[76][152],
reservoir_weight[76][153],
reservoir_weight[76][154],
reservoir_weight[76][155],
reservoir_weight[76][156],
reservoir_weight[76][157],
reservoir_weight[76][158],
reservoir_weight[76][159],
reservoir_weight[76][160],
reservoir_weight[76][161],
reservoir_weight[76][162],
reservoir_weight[76][163],
reservoir_weight[76][164],
reservoir_weight[76][165],
reservoir_weight[76][166],
reservoir_weight[76][167],
reservoir_weight[76][168],
reservoir_weight[76][169],
reservoir_weight[76][170],
reservoir_weight[76][171],
reservoir_weight[76][172],
reservoir_weight[76][173],
reservoir_weight[76][174],
reservoir_weight[76][175],
reservoir_weight[76][176],
reservoir_weight[76][177],
reservoir_weight[76][178],
reservoir_weight[76][179],
reservoir_weight[76][180],
reservoir_weight[76][181],
reservoir_weight[76][182],
reservoir_weight[76][183],
reservoir_weight[76][184],
reservoir_weight[76][185],
reservoir_weight[76][186],
reservoir_weight[76][187],
reservoir_weight[76][188],
reservoir_weight[76][189],
reservoir_weight[76][190],
reservoir_weight[76][191],
reservoir_weight[76][192],
reservoir_weight[76][193],
reservoir_weight[76][194],
reservoir_weight[76][195],
reservoir_weight[76][196],
reservoir_weight[76][197],
reservoir_weight[76][198],
reservoir_weight[76][199]
},
{reservoir_weight[77][0],
reservoir_weight[77][1],
reservoir_weight[77][2],
reservoir_weight[77][3],
reservoir_weight[77][4],
reservoir_weight[77][5],
reservoir_weight[77][6],
reservoir_weight[77][7],
reservoir_weight[77][8],
reservoir_weight[77][9],
reservoir_weight[77][10],
reservoir_weight[77][11],
reservoir_weight[77][12],
reservoir_weight[77][13],
reservoir_weight[77][14],
reservoir_weight[77][15],
reservoir_weight[77][16],
reservoir_weight[77][17],
reservoir_weight[77][18],
reservoir_weight[77][19],
reservoir_weight[77][20],
reservoir_weight[77][21],
reservoir_weight[77][22],
reservoir_weight[77][23],
reservoir_weight[77][24],
reservoir_weight[77][25],
reservoir_weight[77][26],
reservoir_weight[77][27],
reservoir_weight[77][28],
reservoir_weight[77][29],
reservoir_weight[77][30],
reservoir_weight[77][31],
reservoir_weight[77][32],
reservoir_weight[77][33],
reservoir_weight[77][34],
reservoir_weight[77][35],
reservoir_weight[77][36],
reservoir_weight[77][37],
reservoir_weight[77][38],
reservoir_weight[77][39],
reservoir_weight[77][40],
reservoir_weight[77][41],
reservoir_weight[77][42],
reservoir_weight[77][43],
reservoir_weight[77][44],
reservoir_weight[77][45],
reservoir_weight[77][46],
reservoir_weight[77][47],
reservoir_weight[77][48],
reservoir_weight[77][49],
reservoir_weight[77][50],
reservoir_weight[77][51],
reservoir_weight[77][52],
reservoir_weight[77][53],
reservoir_weight[77][54],
reservoir_weight[77][55],
reservoir_weight[77][56],
reservoir_weight[77][57],
reservoir_weight[77][58],
reservoir_weight[77][59],
reservoir_weight[77][60],
reservoir_weight[77][61],
reservoir_weight[77][62],
reservoir_weight[77][63],
reservoir_weight[77][64],
reservoir_weight[77][65],
reservoir_weight[77][66],
reservoir_weight[77][67],
reservoir_weight[77][68],
reservoir_weight[77][69],
reservoir_weight[77][70],
reservoir_weight[77][71],
reservoir_weight[77][72],
reservoir_weight[77][73],
reservoir_weight[77][74],
reservoir_weight[77][75],
reservoir_weight[77][76],
reservoir_weight[77][77],
reservoir_weight[77][78],
reservoir_weight[77][79],
reservoir_weight[77][80],
reservoir_weight[77][81],
reservoir_weight[77][82],
reservoir_weight[77][83],
reservoir_weight[77][84],
reservoir_weight[77][85],
reservoir_weight[77][86],
reservoir_weight[77][87],
reservoir_weight[77][88],
reservoir_weight[77][89],
reservoir_weight[77][90],
reservoir_weight[77][91],
reservoir_weight[77][92],
reservoir_weight[77][93],
reservoir_weight[77][94],
reservoir_weight[77][95],
reservoir_weight[77][96],
reservoir_weight[77][97],
reservoir_weight[77][98],
reservoir_weight[77][99],
reservoir_weight[77][100],
reservoir_weight[77][101],
reservoir_weight[77][102],
reservoir_weight[77][103],
reservoir_weight[77][104],
reservoir_weight[77][105],
reservoir_weight[77][106],
reservoir_weight[77][107],
reservoir_weight[77][108],
reservoir_weight[77][109],
reservoir_weight[77][110],
reservoir_weight[77][111],
reservoir_weight[77][112],
reservoir_weight[77][113],
reservoir_weight[77][114],
reservoir_weight[77][115],
reservoir_weight[77][116],
reservoir_weight[77][117],
reservoir_weight[77][118],
reservoir_weight[77][119],
reservoir_weight[77][120],
reservoir_weight[77][121],
reservoir_weight[77][122],
reservoir_weight[77][123],
reservoir_weight[77][124],
reservoir_weight[77][125],
reservoir_weight[77][126],
reservoir_weight[77][127],
reservoir_weight[77][128],
reservoir_weight[77][129],
reservoir_weight[77][130],
reservoir_weight[77][131],
reservoir_weight[77][132],
reservoir_weight[77][133],
reservoir_weight[77][134],
reservoir_weight[77][135],
reservoir_weight[77][136],
reservoir_weight[77][137],
reservoir_weight[77][138],
reservoir_weight[77][139],
reservoir_weight[77][140],
reservoir_weight[77][141],
reservoir_weight[77][142],
reservoir_weight[77][143],
reservoir_weight[77][144],
reservoir_weight[77][145],
reservoir_weight[77][146],
reservoir_weight[77][147],
reservoir_weight[77][148],
reservoir_weight[77][149],
reservoir_weight[77][150],
reservoir_weight[77][151],
reservoir_weight[77][152],
reservoir_weight[77][153],
reservoir_weight[77][154],
reservoir_weight[77][155],
reservoir_weight[77][156],
reservoir_weight[77][157],
reservoir_weight[77][158],
reservoir_weight[77][159],
reservoir_weight[77][160],
reservoir_weight[77][161],
reservoir_weight[77][162],
reservoir_weight[77][163],
reservoir_weight[77][164],
reservoir_weight[77][165],
reservoir_weight[77][166],
reservoir_weight[77][167],
reservoir_weight[77][168],
reservoir_weight[77][169],
reservoir_weight[77][170],
reservoir_weight[77][171],
reservoir_weight[77][172],
reservoir_weight[77][173],
reservoir_weight[77][174],
reservoir_weight[77][175],
reservoir_weight[77][176],
reservoir_weight[77][177],
reservoir_weight[77][178],
reservoir_weight[77][179],
reservoir_weight[77][180],
reservoir_weight[77][181],
reservoir_weight[77][182],
reservoir_weight[77][183],
reservoir_weight[77][184],
reservoir_weight[77][185],
reservoir_weight[77][186],
reservoir_weight[77][187],
reservoir_weight[77][188],
reservoir_weight[77][189],
reservoir_weight[77][190],
reservoir_weight[77][191],
reservoir_weight[77][192],
reservoir_weight[77][193],
reservoir_weight[77][194],
reservoir_weight[77][195],
reservoir_weight[77][196],
reservoir_weight[77][197],
reservoir_weight[77][198],
reservoir_weight[77][199]
},
{reservoir_weight[78][0],
reservoir_weight[78][1],
reservoir_weight[78][2],
reservoir_weight[78][3],
reservoir_weight[78][4],
reservoir_weight[78][5],
reservoir_weight[78][6],
reservoir_weight[78][7],
reservoir_weight[78][8],
reservoir_weight[78][9],
reservoir_weight[78][10],
reservoir_weight[78][11],
reservoir_weight[78][12],
reservoir_weight[78][13],
reservoir_weight[78][14],
reservoir_weight[78][15],
reservoir_weight[78][16],
reservoir_weight[78][17],
reservoir_weight[78][18],
reservoir_weight[78][19],
reservoir_weight[78][20],
reservoir_weight[78][21],
reservoir_weight[78][22],
reservoir_weight[78][23],
reservoir_weight[78][24],
reservoir_weight[78][25],
reservoir_weight[78][26],
reservoir_weight[78][27],
reservoir_weight[78][28],
reservoir_weight[78][29],
reservoir_weight[78][30],
reservoir_weight[78][31],
reservoir_weight[78][32],
reservoir_weight[78][33],
reservoir_weight[78][34],
reservoir_weight[78][35],
reservoir_weight[78][36],
reservoir_weight[78][37],
reservoir_weight[78][38],
reservoir_weight[78][39],
reservoir_weight[78][40],
reservoir_weight[78][41],
reservoir_weight[78][42],
reservoir_weight[78][43],
reservoir_weight[78][44],
reservoir_weight[78][45],
reservoir_weight[78][46],
reservoir_weight[78][47],
reservoir_weight[78][48],
reservoir_weight[78][49],
reservoir_weight[78][50],
reservoir_weight[78][51],
reservoir_weight[78][52],
reservoir_weight[78][53],
reservoir_weight[78][54],
reservoir_weight[78][55],
reservoir_weight[78][56],
reservoir_weight[78][57],
reservoir_weight[78][58],
reservoir_weight[78][59],
reservoir_weight[78][60],
reservoir_weight[78][61],
reservoir_weight[78][62],
reservoir_weight[78][63],
reservoir_weight[78][64],
reservoir_weight[78][65],
reservoir_weight[78][66],
reservoir_weight[78][67],
reservoir_weight[78][68],
reservoir_weight[78][69],
reservoir_weight[78][70],
reservoir_weight[78][71],
reservoir_weight[78][72],
reservoir_weight[78][73],
reservoir_weight[78][74],
reservoir_weight[78][75],
reservoir_weight[78][76],
reservoir_weight[78][77],
reservoir_weight[78][78],
reservoir_weight[78][79],
reservoir_weight[78][80],
reservoir_weight[78][81],
reservoir_weight[78][82],
reservoir_weight[78][83],
reservoir_weight[78][84],
reservoir_weight[78][85],
reservoir_weight[78][86],
reservoir_weight[78][87],
reservoir_weight[78][88],
reservoir_weight[78][89],
reservoir_weight[78][90],
reservoir_weight[78][91],
reservoir_weight[78][92],
reservoir_weight[78][93],
reservoir_weight[78][94],
reservoir_weight[78][95],
reservoir_weight[78][96],
reservoir_weight[78][97],
reservoir_weight[78][98],
reservoir_weight[78][99],
reservoir_weight[78][100],
reservoir_weight[78][101],
reservoir_weight[78][102],
reservoir_weight[78][103],
reservoir_weight[78][104],
reservoir_weight[78][105],
reservoir_weight[78][106],
reservoir_weight[78][107],
reservoir_weight[78][108],
reservoir_weight[78][109],
reservoir_weight[78][110],
reservoir_weight[78][111],
reservoir_weight[78][112],
reservoir_weight[78][113],
reservoir_weight[78][114],
reservoir_weight[78][115],
reservoir_weight[78][116],
reservoir_weight[78][117],
reservoir_weight[78][118],
reservoir_weight[78][119],
reservoir_weight[78][120],
reservoir_weight[78][121],
reservoir_weight[78][122],
reservoir_weight[78][123],
reservoir_weight[78][124],
reservoir_weight[78][125],
reservoir_weight[78][126],
reservoir_weight[78][127],
reservoir_weight[78][128],
reservoir_weight[78][129],
reservoir_weight[78][130],
reservoir_weight[78][131],
reservoir_weight[78][132],
reservoir_weight[78][133],
reservoir_weight[78][134],
reservoir_weight[78][135],
reservoir_weight[78][136],
reservoir_weight[78][137],
reservoir_weight[78][138],
reservoir_weight[78][139],
reservoir_weight[78][140],
reservoir_weight[78][141],
reservoir_weight[78][142],
reservoir_weight[78][143],
reservoir_weight[78][144],
reservoir_weight[78][145],
reservoir_weight[78][146],
reservoir_weight[78][147],
reservoir_weight[78][148],
reservoir_weight[78][149],
reservoir_weight[78][150],
reservoir_weight[78][151],
reservoir_weight[78][152],
reservoir_weight[78][153],
reservoir_weight[78][154],
reservoir_weight[78][155],
reservoir_weight[78][156],
reservoir_weight[78][157],
reservoir_weight[78][158],
reservoir_weight[78][159],
reservoir_weight[78][160],
reservoir_weight[78][161],
reservoir_weight[78][162],
reservoir_weight[78][163],
reservoir_weight[78][164],
reservoir_weight[78][165],
reservoir_weight[78][166],
reservoir_weight[78][167],
reservoir_weight[78][168],
reservoir_weight[78][169],
reservoir_weight[78][170],
reservoir_weight[78][171],
reservoir_weight[78][172],
reservoir_weight[78][173],
reservoir_weight[78][174],
reservoir_weight[78][175],
reservoir_weight[78][176],
reservoir_weight[78][177],
reservoir_weight[78][178],
reservoir_weight[78][179],
reservoir_weight[78][180],
reservoir_weight[78][181],
reservoir_weight[78][182],
reservoir_weight[78][183],
reservoir_weight[78][184],
reservoir_weight[78][185],
reservoir_weight[78][186],
reservoir_weight[78][187],
reservoir_weight[78][188],
reservoir_weight[78][189],
reservoir_weight[78][190],
reservoir_weight[78][191],
reservoir_weight[78][192],
reservoir_weight[78][193],
reservoir_weight[78][194],
reservoir_weight[78][195],
reservoir_weight[78][196],
reservoir_weight[78][197],
reservoir_weight[78][198],
reservoir_weight[78][199]
},
{reservoir_weight[79][0],
reservoir_weight[79][1],
reservoir_weight[79][2],
reservoir_weight[79][3],
reservoir_weight[79][4],
reservoir_weight[79][5],
reservoir_weight[79][6],
reservoir_weight[79][7],
reservoir_weight[79][8],
reservoir_weight[79][9],
reservoir_weight[79][10],
reservoir_weight[79][11],
reservoir_weight[79][12],
reservoir_weight[79][13],
reservoir_weight[79][14],
reservoir_weight[79][15],
reservoir_weight[79][16],
reservoir_weight[79][17],
reservoir_weight[79][18],
reservoir_weight[79][19],
reservoir_weight[79][20],
reservoir_weight[79][21],
reservoir_weight[79][22],
reservoir_weight[79][23],
reservoir_weight[79][24],
reservoir_weight[79][25],
reservoir_weight[79][26],
reservoir_weight[79][27],
reservoir_weight[79][28],
reservoir_weight[79][29],
reservoir_weight[79][30],
reservoir_weight[79][31],
reservoir_weight[79][32],
reservoir_weight[79][33],
reservoir_weight[79][34],
reservoir_weight[79][35],
reservoir_weight[79][36],
reservoir_weight[79][37],
reservoir_weight[79][38],
reservoir_weight[79][39],
reservoir_weight[79][40],
reservoir_weight[79][41],
reservoir_weight[79][42],
reservoir_weight[79][43],
reservoir_weight[79][44],
reservoir_weight[79][45],
reservoir_weight[79][46],
reservoir_weight[79][47],
reservoir_weight[79][48],
reservoir_weight[79][49],
reservoir_weight[79][50],
reservoir_weight[79][51],
reservoir_weight[79][52],
reservoir_weight[79][53],
reservoir_weight[79][54],
reservoir_weight[79][55],
reservoir_weight[79][56],
reservoir_weight[79][57],
reservoir_weight[79][58],
reservoir_weight[79][59],
reservoir_weight[79][60],
reservoir_weight[79][61],
reservoir_weight[79][62],
reservoir_weight[79][63],
reservoir_weight[79][64],
reservoir_weight[79][65],
reservoir_weight[79][66],
reservoir_weight[79][67],
reservoir_weight[79][68],
reservoir_weight[79][69],
reservoir_weight[79][70],
reservoir_weight[79][71],
reservoir_weight[79][72],
reservoir_weight[79][73],
reservoir_weight[79][74],
reservoir_weight[79][75],
reservoir_weight[79][76],
reservoir_weight[79][77],
reservoir_weight[79][78],
reservoir_weight[79][79],
reservoir_weight[79][80],
reservoir_weight[79][81],
reservoir_weight[79][82],
reservoir_weight[79][83],
reservoir_weight[79][84],
reservoir_weight[79][85],
reservoir_weight[79][86],
reservoir_weight[79][87],
reservoir_weight[79][88],
reservoir_weight[79][89],
reservoir_weight[79][90],
reservoir_weight[79][91],
reservoir_weight[79][92],
reservoir_weight[79][93],
reservoir_weight[79][94],
reservoir_weight[79][95],
reservoir_weight[79][96],
reservoir_weight[79][97],
reservoir_weight[79][98],
reservoir_weight[79][99],
reservoir_weight[79][100],
reservoir_weight[79][101],
reservoir_weight[79][102],
reservoir_weight[79][103],
reservoir_weight[79][104],
reservoir_weight[79][105],
reservoir_weight[79][106],
reservoir_weight[79][107],
reservoir_weight[79][108],
reservoir_weight[79][109],
reservoir_weight[79][110],
reservoir_weight[79][111],
reservoir_weight[79][112],
reservoir_weight[79][113],
reservoir_weight[79][114],
reservoir_weight[79][115],
reservoir_weight[79][116],
reservoir_weight[79][117],
reservoir_weight[79][118],
reservoir_weight[79][119],
reservoir_weight[79][120],
reservoir_weight[79][121],
reservoir_weight[79][122],
reservoir_weight[79][123],
reservoir_weight[79][124],
reservoir_weight[79][125],
reservoir_weight[79][126],
reservoir_weight[79][127],
reservoir_weight[79][128],
reservoir_weight[79][129],
reservoir_weight[79][130],
reservoir_weight[79][131],
reservoir_weight[79][132],
reservoir_weight[79][133],
reservoir_weight[79][134],
reservoir_weight[79][135],
reservoir_weight[79][136],
reservoir_weight[79][137],
reservoir_weight[79][138],
reservoir_weight[79][139],
reservoir_weight[79][140],
reservoir_weight[79][141],
reservoir_weight[79][142],
reservoir_weight[79][143],
reservoir_weight[79][144],
reservoir_weight[79][145],
reservoir_weight[79][146],
reservoir_weight[79][147],
reservoir_weight[79][148],
reservoir_weight[79][149],
reservoir_weight[79][150],
reservoir_weight[79][151],
reservoir_weight[79][152],
reservoir_weight[79][153],
reservoir_weight[79][154],
reservoir_weight[79][155],
reservoir_weight[79][156],
reservoir_weight[79][157],
reservoir_weight[79][158],
reservoir_weight[79][159],
reservoir_weight[79][160],
reservoir_weight[79][161],
reservoir_weight[79][162],
reservoir_weight[79][163],
reservoir_weight[79][164],
reservoir_weight[79][165],
reservoir_weight[79][166],
reservoir_weight[79][167],
reservoir_weight[79][168],
reservoir_weight[79][169],
reservoir_weight[79][170],
reservoir_weight[79][171],
reservoir_weight[79][172],
reservoir_weight[79][173],
reservoir_weight[79][174],
reservoir_weight[79][175],
reservoir_weight[79][176],
reservoir_weight[79][177],
reservoir_weight[79][178],
reservoir_weight[79][179],
reservoir_weight[79][180],
reservoir_weight[79][181],
reservoir_weight[79][182],
reservoir_weight[79][183],
reservoir_weight[79][184],
reservoir_weight[79][185],
reservoir_weight[79][186],
reservoir_weight[79][187],
reservoir_weight[79][188],
reservoir_weight[79][189],
reservoir_weight[79][190],
reservoir_weight[79][191],
reservoir_weight[79][192],
reservoir_weight[79][193],
reservoir_weight[79][194],
reservoir_weight[79][195],
reservoir_weight[79][196],
reservoir_weight[79][197],
reservoir_weight[79][198],
reservoir_weight[79][199]
},
{reservoir_weight[80][0],
reservoir_weight[80][1],
reservoir_weight[80][2],
reservoir_weight[80][3],
reservoir_weight[80][4],
reservoir_weight[80][5],
reservoir_weight[80][6],
reservoir_weight[80][7],
reservoir_weight[80][8],
reservoir_weight[80][9],
reservoir_weight[80][10],
reservoir_weight[80][11],
reservoir_weight[80][12],
reservoir_weight[80][13],
reservoir_weight[80][14],
reservoir_weight[80][15],
reservoir_weight[80][16],
reservoir_weight[80][17],
reservoir_weight[80][18],
reservoir_weight[80][19],
reservoir_weight[80][20],
reservoir_weight[80][21],
reservoir_weight[80][22],
reservoir_weight[80][23],
reservoir_weight[80][24],
reservoir_weight[80][25],
reservoir_weight[80][26],
reservoir_weight[80][27],
reservoir_weight[80][28],
reservoir_weight[80][29],
reservoir_weight[80][30],
reservoir_weight[80][31],
reservoir_weight[80][32],
reservoir_weight[80][33],
reservoir_weight[80][34],
reservoir_weight[80][35],
reservoir_weight[80][36],
reservoir_weight[80][37],
reservoir_weight[80][38],
reservoir_weight[80][39],
reservoir_weight[80][40],
reservoir_weight[80][41],
reservoir_weight[80][42],
reservoir_weight[80][43],
reservoir_weight[80][44],
reservoir_weight[80][45],
reservoir_weight[80][46],
reservoir_weight[80][47],
reservoir_weight[80][48],
reservoir_weight[80][49],
reservoir_weight[80][50],
reservoir_weight[80][51],
reservoir_weight[80][52],
reservoir_weight[80][53],
reservoir_weight[80][54],
reservoir_weight[80][55],
reservoir_weight[80][56],
reservoir_weight[80][57],
reservoir_weight[80][58],
reservoir_weight[80][59],
reservoir_weight[80][60],
reservoir_weight[80][61],
reservoir_weight[80][62],
reservoir_weight[80][63],
reservoir_weight[80][64],
reservoir_weight[80][65],
reservoir_weight[80][66],
reservoir_weight[80][67],
reservoir_weight[80][68],
reservoir_weight[80][69],
reservoir_weight[80][70],
reservoir_weight[80][71],
reservoir_weight[80][72],
reservoir_weight[80][73],
reservoir_weight[80][74],
reservoir_weight[80][75],
reservoir_weight[80][76],
reservoir_weight[80][77],
reservoir_weight[80][78],
reservoir_weight[80][79],
reservoir_weight[80][80],
reservoir_weight[80][81],
reservoir_weight[80][82],
reservoir_weight[80][83],
reservoir_weight[80][84],
reservoir_weight[80][85],
reservoir_weight[80][86],
reservoir_weight[80][87],
reservoir_weight[80][88],
reservoir_weight[80][89],
reservoir_weight[80][90],
reservoir_weight[80][91],
reservoir_weight[80][92],
reservoir_weight[80][93],
reservoir_weight[80][94],
reservoir_weight[80][95],
reservoir_weight[80][96],
reservoir_weight[80][97],
reservoir_weight[80][98],
reservoir_weight[80][99],
reservoir_weight[80][100],
reservoir_weight[80][101],
reservoir_weight[80][102],
reservoir_weight[80][103],
reservoir_weight[80][104],
reservoir_weight[80][105],
reservoir_weight[80][106],
reservoir_weight[80][107],
reservoir_weight[80][108],
reservoir_weight[80][109],
reservoir_weight[80][110],
reservoir_weight[80][111],
reservoir_weight[80][112],
reservoir_weight[80][113],
reservoir_weight[80][114],
reservoir_weight[80][115],
reservoir_weight[80][116],
reservoir_weight[80][117],
reservoir_weight[80][118],
reservoir_weight[80][119],
reservoir_weight[80][120],
reservoir_weight[80][121],
reservoir_weight[80][122],
reservoir_weight[80][123],
reservoir_weight[80][124],
reservoir_weight[80][125],
reservoir_weight[80][126],
reservoir_weight[80][127],
reservoir_weight[80][128],
reservoir_weight[80][129],
reservoir_weight[80][130],
reservoir_weight[80][131],
reservoir_weight[80][132],
reservoir_weight[80][133],
reservoir_weight[80][134],
reservoir_weight[80][135],
reservoir_weight[80][136],
reservoir_weight[80][137],
reservoir_weight[80][138],
reservoir_weight[80][139],
reservoir_weight[80][140],
reservoir_weight[80][141],
reservoir_weight[80][142],
reservoir_weight[80][143],
reservoir_weight[80][144],
reservoir_weight[80][145],
reservoir_weight[80][146],
reservoir_weight[80][147],
reservoir_weight[80][148],
reservoir_weight[80][149],
reservoir_weight[80][150],
reservoir_weight[80][151],
reservoir_weight[80][152],
reservoir_weight[80][153],
reservoir_weight[80][154],
reservoir_weight[80][155],
reservoir_weight[80][156],
reservoir_weight[80][157],
reservoir_weight[80][158],
reservoir_weight[80][159],
reservoir_weight[80][160],
reservoir_weight[80][161],
reservoir_weight[80][162],
reservoir_weight[80][163],
reservoir_weight[80][164],
reservoir_weight[80][165],
reservoir_weight[80][166],
reservoir_weight[80][167],
reservoir_weight[80][168],
reservoir_weight[80][169],
reservoir_weight[80][170],
reservoir_weight[80][171],
reservoir_weight[80][172],
reservoir_weight[80][173],
reservoir_weight[80][174],
reservoir_weight[80][175],
reservoir_weight[80][176],
reservoir_weight[80][177],
reservoir_weight[80][178],
reservoir_weight[80][179],
reservoir_weight[80][180],
reservoir_weight[80][181],
reservoir_weight[80][182],
reservoir_weight[80][183],
reservoir_weight[80][184],
reservoir_weight[80][185],
reservoir_weight[80][186],
reservoir_weight[80][187],
reservoir_weight[80][188],
reservoir_weight[80][189],
reservoir_weight[80][190],
reservoir_weight[80][191],
reservoir_weight[80][192],
reservoir_weight[80][193],
reservoir_weight[80][194],
reservoir_weight[80][195],
reservoir_weight[80][196],
reservoir_weight[80][197],
reservoir_weight[80][198],
reservoir_weight[80][199]
},
{reservoir_weight[81][0],
reservoir_weight[81][1],
reservoir_weight[81][2],
reservoir_weight[81][3],
reservoir_weight[81][4],
reservoir_weight[81][5],
reservoir_weight[81][6],
reservoir_weight[81][7],
reservoir_weight[81][8],
reservoir_weight[81][9],
reservoir_weight[81][10],
reservoir_weight[81][11],
reservoir_weight[81][12],
reservoir_weight[81][13],
reservoir_weight[81][14],
reservoir_weight[81][15],
reservoir_weight[81][16],
reservoir_weight[81][17],
reservoir_weight[81][18],
reservoir_weight[81][19],
reservoir_weight[81][20],
reservoir_weight[81][21],
reservoir_weight[81][22],
reservoir_weight[81][23],
reservoir_weight[81][24],
reservoir_weight[81][25],
reservoir_weight[81][26],
reservoir_weight[81][27],
reservoir_weight[81][28],
reservoir_weight[81][29],
reservoir_weight[81][30],
reservoir_weight[81][31],
reservoir_weight[81][32],
reservoir_weight[81][33],
reservoir_weight[81][34],
reservoir_weight[81][35],
reservoir_weight[81][36],
reservoir_weight[81][37],
reservoir_weight[81][38],
reservoir_weight[81][39],
reservoir_weight[81][40],
reservoir_weight[81][41],
reservoir_weight[81][42],
reservoir_weight[81][43],
reservoir_weight[81][44],
reservoir_weight[81][45],
reservoir_weight[81][46],
reservoir_weight[81][47],
reservoir_weight[81][48],
reservoir_weight[81][49],
reservoir_weight[81][50],
reservoir_weight[81][51],
reservoir_weight[81][52],
reservoir_weight[81][53],
reservoir_weight[81][54],
reservoir_weight[81][55],
reservoir_weight[81][56],
reservoir_weight[81][57],
reservoir_weight[81][58],
reservoir_weight[81][59],
reservoir_weight[81][60],
reservoir_weight[81][61],
reservoir_weight[81][62],
reservoir_weight[81][63],
reservoir_weight[81][64],
reservoir_weight[81][65],
reservoir_weight[81][66],
reservoir_weight[81][67],
reservoir_weight[81][68],
reservoir_weight[81][69],
reservoir_weight[81][70],
reservoir_weight[81][71],
reservoir_weight[81][72],
reservoir_weight[81][73],
reservoir_weight[81][74],
reservoir_weight[81][75],
reservoir_weight[81][76],
reservoir_weight[81][77],
reservoir_weight[81][78],
reservoir_weight[81][79],
reservoir_weight[81][80],
reservoir_weight[81][81],
reservoir_weight[81][82],
reservoir_weight[81][83],
reservoir_weight[81][84],
reservoir_weight[81][85],
reservoir_weight[81][86],
reservoir_weight[81][87],
reservoir_weight[81][88],
reservoir_weight[81][89],
reservoir_weight[81][90],
reservoir_weight[81][91],
reservoir_weight[81][92],
reservoir_weight[81][93],
reservoir_weight[81][94],
reservoir_weight[81][95],
reservoir_weight[81][96],
reservoir_weight[81][97],
reservoir_weight[81][98],
reservoir_weight[81][99],
reservoir_weight[81][100],
reservoir_weight[81][101],
reservoir_weight[81][102],
reservoir_weight[81][103],
reservoir_weight[81][104],
reservoir_weight[81][105],
reservoir_weight[81][106],
reservoir_weight[81][107],
reservoir_weight[81][108],
reservoir_weight[81][109],
reservoir_weight[81][110],
reservoir_weight[81][111],
reservoir_weight[81][112],
reservoir_weight[81][113],
reservoir_weight[81][114],
reservoir_weight[81][115],
reservoir_weight[81][116],
reservoir_weight[81][117],
reservoir_weight[81][118],
reservoir_weight[81][119],
reservoir_weight[81][120],
reservoir_weight[81][121],
reservoir_weight[81][122],
reservoir_weight[81][123],
reservoir_weight[81][124],
reservoir_weight[81][125],
reservoir_weight[81][126],
reservoir_weight[81][127],
reservoir_weight[81][128],
reservoir_weight[81][129],
reservoir_weight[81][130],
reservoir_weight[81][131],
reservoir_weight[81][132],
reservoir_weight[81][133],
reservoir_weight[81][134],
reservoir_weight[81][135],
reservoir_weight[81][136],
reservoir_weight[81][137],
reservoir_weight[81][138],
reservoir_weight[81][139],
reservoir_weight[81][140],
reservoir_weight[81][141],
reservoir_weight[81][142],
reservoir_weight[81][143],
reservoir_weight[81][144],
reservoir_weight[81][145],
reservoir_weight[81][146],
reservoir_weight[81][147],
reservoir_weight[81][148],
reservoir_weight[81][149],
reservoir_weight[81][150],
reservoir_weight[81][151],
reservoir_weight[81][152],
reservoir_weight[81][153],
reservoir_weight[81][154],
reservoir_weight[81][155],
reservoir_weight[81][156],
reservoir_weight[81][157],
reservoir_weight[81][158],
reservoir_weight[81][159],
reservoir_weight[81][160],
reservoir_weight[81][161],
reservoir_weight[81][162],
reservoir_weight[81][163],
reservoir_weight[81][164],
reservoir_weight[81][165],
reservoir_weight[81][166],
reservoir_weight[81][167],
reservoir_weight[81][168],
reservoir_weight[81][169],
reservoir_weight[81][170],
reservoir_weight[81][171],
reservoir_weight[81][172],
reservoir_weight[81][173],
reservoir_weight[81][174],
reservoir_weight[81][175],
reservoir_weight[81][176],
reservoir_weight[81][177],
reservoir_weight[81][178],
reservoir_weight[81][179],
reservoir_weight[81][180],
reservoir_weight[81][181],
reservoir_weight[81][182],
reservoir_weight[81][183],
reservoir_weight[81][184],
reservoir_weight[81][185],
reservoir_weight[81][186],
reservoir_weight[81][187],
reservoir_weight[81][188],
reservoir_weight[81][189],
reservoir_weight[81][190],
reservoir_weight[81][191],
reservoir_weight[81][192],
reservoir_weight[81][193],
reservoir_weight[81][194],
reservoir_weight[81][195],
reservoir_weight[81][196],
reservoir_weight[81][197],
reservoir_weight[81][198],
reservoir_weight[81][199]
},
{reservoir_weight[82][0],
reservoir_weight[82][1],
reservoir_weight[82][2],
reservoir_weight[82][3],
reservoir_weight[82][4],
reservoir_weight[82][5],
reservoir_weight[82][6],
reservoir_weight[82][7],
reservoir_weight[82][8],
reservoir_weight[82][9],
reservoir_weight[82][10],
reservoir_weight[82][11],
reservoir_weight[82][12],
reservoir_weight[82][13],
reservoir_weight[82][14],
reservoir_weight[82][15],
reservoir_weight[82][16],
reservoir_weight[82][17],
reservoir_weight[82][18],
reservoir_weight[82][19],
reservoir_weight[82][20],
reservoir_weight[82][21],
reservoir_weight[82][22],
reservoir_weight[82][23],
reservoir_weight[82][24],
reservoir_weight[82][25],
reservoir_weight[82][26],
reservoir_weight[82][27],
reservoir_weight[82][28],
reservoir_weight[82][29],
reservoir_weight[82][30],
reservoir_weight[82][31],
reservoir_weight[82][32],
reservoir_weight[82][33],
reservoir_weight[82][34],
reservoir_weight[82][35],
reservoir_weight[82][36],
reservoir_weight[82][37],
reservoir_weight[82][38],
reservoir_weight[82][39],
reservoir_weight[82][40],
reservoir_weight[82][41],
reservoir_weight[82][42],
reservoir_weight[82][43],
reservoir_weight[82][44],
reservoir_weight[82][45],
reservoir_weight[82][46],
reservoir_weight[82][47],
reservoir_weight[82][48],
reservoir_weight[82][49],
reservoir_weight[82][50],
reservoir_weight[82][51],
reservoir_weight[82][52],
reservoir_weight[82][53],
reservoir_weight[82][54],
reservoir_weight[82][55],
reservoir_weight[82][56],
reservoir_weight[82][57],
reservoir_weight[82][58],
reservoir_weight[82][59],
reservoir_weight[82][60],
reservoir_weight[82][61],
reservoir_weight[82][62],
reservoir_weight[82][63],
reservoir_weight[82][64],
reservoir_weight[82][65],
reservoir_weight[82][66],
reservoir_weight[82][67],
reservoir_weight[82][68],
reservoir_weight[82][69],
reservoir_weight[82][70],
reservoir_weight[82][71],
reservoir_weight[82][72],
reservoir_weight[82][73],
reservoir_weight[82][74],
reservoir_weight[82][75],
reservoir_weight[82][76],
reservoir_weight[82][77],
reservoir_weight[82][78],
reservoir_weight[82][79],
reservoir_weight[82][80],
reservoir_weight[82][81],
reservoir_weight[82][82],
reservoir_weight[82][83],
reservoir_weight[82][84],
reservoir_weight[82][85],
reservoir_weight[82][86],
reservoir_weight[82][87],
reservoir_weight[82][88],
reservoir_weight[82][89],
reservoir_weight[82][90],
reservoir_weight[82][91],
reservoir_weight[82][92],
reservoir_weight[82][93],
reservoir_weight[82][94],
reservoir_weight[82][95],
reservoir_weight[82][96],
reservoir_weight[82][97],
reservoir_weight[82][98],
reservoir_weight[82][99],
reservoir_weight[82][100],
reservoir_weight[82][101],
reservoir_weight[82][102],
reservoir_weight[82][103],
reservoir_weight[82][104],
reservoir_weight[82][105],
reservoir_weight[82][106],
reservoir_weight[82][107],
reservoir_weight[82][108],
reservoir_weight[82][109],
reservoir_weight[82][110],
reservoir_weight[82][111],
reservoir_weight[82][112],
reservoir_weight[82][113],
reservoir_weight[82][114],
reservoir_weight[82][115],
reservoir_weight[82][116],
reservoir_weight[82][117],
reservoir_weight[82][118],
reservoir_weight[82][119],
reservoir_weight[82][120],
reservoir_weight[82][121],
reservoir_weight[82][122],
reservoir_weight[82][123],
reservoir_weight[82][124],
reservoir_weight[82][125],
reservoir_weight[82][126],
reservoir_weight[82][127],
reservoir_weight[82][128],
reservoir_weight[82][129],
reservoir_weight[82][130],
reservoir_weight[82][131],
reservoir_weight[82][132],
reservoir_weight[82][133],
reservoir_weight[82][134],
reservoir_weight[82][135],
reservoir_weight[82][136],
reservoir_weight[82][137],
reservoir_weight[82][138],
reservoir_weight[82][139],
reservoir_weight[82][140],
reservoir_weight[82][141],
reservoir_weight[82][142],
reservoir_weight[82][143],
reservoir_weight[82][144],
reservoir_weight[82][145],
reservoir_weight[82][146],
reservoir_weight[82][147],
reservoir_weight[82][148],
reservoir_weight[82][149],
reservoir_weight[82][150],
reservoir_weight[82][151],
reservoir_weight[82][152],
reservoir_weight[82][153],
reservoir_weight[82][154],
reservoir_weight[82][155],
reservoir_weight[82][156],
reservoir_weight[82][157],
reservoir_weight[82][158],
reservoir_weight[82][159],
reservoir_weight[82][160],
reservoir_weight[82][161],
reservoir_weight[82][162],
reservoir_weight[82][163],
reservoir_weight[82][164],
reservoir_weight[82][165],
reservoir_weight[82][166],
reservoir_weight[82][167],
reservoir_weight[82][168],
reservoir_weight[82][169],
reservoir_weight[82][170],
reservoir_weight[82][171],
reservoir_weight[82][172],
reservoir_weight[82][173],
reservoir_weight[82][174],
reservoir_weight[82][175],
reservoir_weight[82][176],
reservoir_weight[82][177],
reservoir_weight[82][178],
reservoir_weight[82][179],
reservoir_weight[82][180],
reservoir_weight[82][181],
reservoir_weight[82][182],
reservoir_weight[82][183],
reservoir_weight[82][184],
reservoir_weight[82][185],
reservoir_weight[82][186],
reservoir_weight[82][187],
reservoir_weight[82][188],
reservoir_weight[82][189],
reservoir_weight[82][190],
reservoir_weight[82][191],
reservoir_weight[82][192],
reservoir_weight[82][193],
reservoir_weight[82][194],
reservoir_weight[82][195],
reservoir_weight[82][196],
reservoir_weight[82][197],
reservoir_weight[82][198],
reservoir_weight[82][199]
},
{reservoir_weight[83][0],
reservoir_weight[83][1],
reservoir_weight[83][2],
reservoir_weight[83][3],
reservoir_weight[83][4],
reservoir_weight[83][5],
reservoir_weight[83][6],
reservoir_weight[83][7],
reservoir_weight[83][8],
reservoir_weight[83][9],
reservoir_weight[83][10],
reservoir_weight[83][11],
reservoir_weight[83][12],
reservoir_weight[83][13],
reservoir_weight[83][14],
reservoir_weight[83][15],
reservoir_weight[83][16],
reservoir_weight[83][17],
reservoir_weight[83][18],
reservoir_weight[83][19],
reservoir_weight[83][20],
reservoir_weight[83][21],
reservoir_weight[83][22],
reservoir_weight[83][23],
reservoir_weight[83][24],
reservoir_weight[83][25],
reservoir_weight[83][26],
reservoir_weight[83][27],
reservoir_weight[83][28],
reservoir_weight[83][29],
reservoir_weight[83][30],
reservoir_weight[83][31],
reservoir_weight[83][32],
reservoir_weight[83][33],
reservoir_weight[83][34],
reservoir_weight[83][35],
reservoir_weight[83][36],
reservoir_weight[83][37],
reservoir_weight[83][38],
reservoir_weight[83][39],
reservoir_weight[83][40],
reservoir_weight[83][41],
reservoir_weight[83][42],
reservoir_weight[83][43],
reservoir_weight[83][44],
reservoir_weight[83][45],
reservoir_weight[83][46],
reservoir_weight[83][47],
reservoir_weight[83][48],
reservoir_weight[83][49],
reservoir_weight[83][50],
reservoir_weight[83][51],
reservoir_weight[83][52],
reservoir_weight[83][53],
reservoir_weight[83][54],
reservoir_weight[83][55],
reservoir_weight[83][56],
reservoir_weight[83][57],
reservoir_weight[83][58],
reservoir_weight[83][59],
reservoir_weight[83][60],
reservoir_weight[83][61],
reservoir_weight[83][62],
reservoir_weight[83][63],
reservoir_weight[83][64],
reservoir_weight[83][65],
reservoir_weight[83][66],
reservoir_weight[83][67],
reservoir_weight[83][68],
reservoir_weight[83][69],
reservoir_weight[83][70],
reservoir_weight[83][71],
reservoir_weight[83][72],
reservoir_weight[83][73],
reservoir_weight[83][74],
reservoir_weight[83][75],
reservoir_weight[83][76],
reservoir_weight[83][77],
reservoir_weight[83][78],
reservoir_weight[83][79],
reservoir_weight[83][80],
reservoir_weight[83][81],
reservoir_weight[83][82],
reservoir_weight[83][83],
reservoir_weight[83][84],
reservoir_weight[83][85],
reservoir_weight[83][86],
reservoir_weight[83][87],
reservoir_weight[83][88],
reservoir_weight[83][89],
reservoir_weight[83][90],
reservoir_weight[83][91],
reservoir_weight[83][92],
reservoir_weight[83][93],
reservoir_weight[83][94],
reservoir_weight[83][95],
reservoir_weight[83][96],
reservoir_weight[83][97],
reservoir_weight[83][98],
reservoir_weight[83][99],
reservoir_weight[83][100],
reservoir_weight[83][101],
reservoir_weight[83][102],
reservoir_weight[83][103],
reservoir_weight[83][104],
reservoir_weight[83][105],
reservoir_weight[83][106],
reservoir_weight[83][107],
reservoir_weight[83][108],
reservoir_weight[83][109],
reservoir_weight[83][110],
reservoir_weight[83][111],
reservoir_weight[83][112],
reservoir_weight[83][113],
reservoir_weight[83][114],
reservoir_weight[83][115],
reservoir_weight[83][116],
reservoir_weight[83][117],
reservoir_weight[83][118],
reservoir_weight[83][119],
reservoir_weight[83][120],
reservoir_weight[83][121],
reservoir_weight[83][122],
reservoir_weight[83][123],
reservoir_weight[83][124],
reservoir_weight[83][125],
reservoir_weight[83][126],
reservoir_weight[83][127],
reservoir_weight[83][128],
reservoir_weight[83][129],
reservoir_weight[83][130],
reservoir_weight[83][131],
reservoir_weight[83][132],
reservoir_weight[83][133],
reservoir_weight[83][134],
reservoir_weight[83][135],
reservoir_weight[83][136],
reservoir_weight[83][137],
reservoir_weight[83][138],
reservoir_weight[83][139],
reservoir_weight[83][140],
reservoir_weight[83][141],
reservoir_weight[83][142],
reservoir_weight[83][143],
reservoir_weight[83][144],
reservoir_weight[83][145],
reservoir_weight[83][146],
reservoir_weight[83][147],
reservoir_weight[83][148],
reservoir_weight[83][149],
reservoir_weight[83][150],
reservoir_weight[83][151],
reservoir_weight[83][152],
reservoir_weight[83][153],
reservoir_weight[83][154],
reservoir_weight[83][155],
reservoir_weight[83][156],
reservoir_weight[83][157],
reservoir_weight[83][158],
reservoir_weight[83][159],
reservoir_weight[83][160],
reservoir_weight[83][161],
reservoir_weight[83][162],
reservoir_weight[83][163],
reservoir_weight[83][164],
reservoir_weight[83][165],
reservoir_weight[83][166],
reservoir_weight[83][167],
reservoir_weight[83][168],
reservoir_weight[83][169],
reservoir_weight[83][170],
reservoir_weight[83][171],
reservoir_weight[83][172],
reservoir_weight[83][173],
reservoir_weight[83][174],
reservoir_weight[83][175],
reservoir_weight[83][176],
reservoir_weight[83][177],
reservoir_weight[83][178],
reservoir_weight[83][179],
reservoir_weight[83][180],
reservoir_weight[83][181],
reservoir_weight[83][182],
reservoir_weight[83][183],
reservoir_weight[83][184],
reservoir_weight[83][185],
reservoir_weight[83][186],
reservoir_weight[83][187],
reservoir_weight[83][188],
reservoir_weight[83][189],
reservoir_weight[83][190],
reservoir_weight[83][191],
reservoir_weight[83][192],
reservoir_weight[83][193],
reservoir_weight[83][194],
reservoir_weight[83][195],
reservoir_weight[83][196],
reservoir_weight[83][197],
reservoir_weight[83][198],
reservoir_weight[83][199]
},
{reservoir_weight[84][0],
reservoir_weight[84][1],
reservoir_weight[84][2],
reservoir_weight[84][3],
reservoir_weight[84][4],
reservoir_weight[84][5],
reservoir_weight[84][6],
reservoir_weight[84][7],
reservoir_weight[84][8],
reservoir_weight[84][9],
reservoir_weight[84][10],
reservoir_weight[84][11],
reservoir_weight[84][12],
reservoir_weight[84][13],
reservoir_weight[84][14],
reservoir_weight[84][15],
reservoir_weight[84][16],
reservoir_weight[84][17],
reservoir_weight[84][18],
reservoir_weight[84][19],
reservoir_weight[84][20],
reservoir_weight[84][21],
reservoir_weight[84][22],
reservoir_weight[84][23],
reservoir_weight[84][24],
reservoir_weight[84][25],
reservoir_weight[84][26],
reservoir_weight[84][27],
reservoir_weight[84][28],
reservoir_weight[84][29],
reservoir_weight[84][30],
reservoir_weight[84][31],
reservoir_weight[84][32],
reservoir_weight[84][33],
reservoir_weight[84][34],
reservoir_weight[84][35],
reservoir_weight[84][36],
reservoir_weight[84][37],
reservoir_weight[84][38],
reservoir_weight[84][39],
reservoir_weight[84][40],
reservoir_weight[84][41],
reservoir_weight[84][42],
reservoir_weight[84][43],
reservoir_weight[84][44],
reservoir_weight[84][45],
reservoir_weight[84][46],
reservoir_weight[84][47],
reservoir_weight[84][48],
reservoir_weight[84][49],
reservoir_weight[84][50],
reservoir_weight[84][51],
reservoir_weight[84][52],
reservoir_weight[84][53],
reservoir_weight[84][54],
reservoir_weight[84][55],
reservoir_weight[84][56],
reservoir_weight[84][57],
reservoir_weight[84][58],
reservoir_weight[84][59],
reservoir_weight[84][60],
reservoir_weight[84][61],
reservoir_weight[84][62],
reservoir_weight[84][63],
reservoir_weight[84][64],
reservoir_weight[84][65],
reservoir_weight[84][66],
reservoir_weight[84][67],
reservoir_weight[84][68],
reservoir_weight[84][69],
reservoir_weight[84][70],
reservoir_weight[84][71],
reservoir_weight[84][72],
reservoir_weight[84][73],
reservoir_weight[84][74],
reservoir_weight[84][75],
reservoir_weight[84][76],
reservoir_weight[84][77],
reservoir_weight[84][78],
reservoir_weight[84][79],
reservoir_weight[84][80],
reservoir_weight[84][81],
reservoir_weight[84][82],
reservoir_weight[84][83],
reservoir_weight[84][84],
reservoir_weight[84][85],
reservoir_weight[84][86],
reservoir_weight[84][87],
reservoir_weight[84][88],
reservoir_weight[84][89],
reservoir_weight[84][90],
reservoir_weight[84][91],
reservoir_weight[84][92],
reservoir_weight[84][93],
reservoir_weight[84][94],
reservoir_weight[84][95],
reservoir_weight[84][96],
reservoir_weight[84][97],
reservoir_weight[84][98],
reservoir_weight[84][99],
reservoir_weight[84][100],
reservoir_weight[84][101],
reservoir_weight[84][102],
reservoir_weight[84][103],
reservoir_weight[84][104],
reservoir_weight[84][105],
reservoir_weight[84][106],
reservoir_weight[84][107],
reservoir_weight[84][108],
reservoir_weight[84][109],
reservoir_weight[84][110],
reservoir_weight[84][111],
reservoir_weight[84][112],
reservoir_weight[84][113],
reservoir_weight[84][114],
reservoir_weight[84][115],
reservoir_weight[84][116],
reservoir_weight[84][117],
reservoir_weight[84][118],
reservoir_weight[84][119],
reservoir_weight[84][120],
reservoir_weight[84][121],
reservoir_weight[84][122],
reservoir_weight[84][123],
reservoir_weight[84][124],
reservoir_weight[84][125],
reservoir_weight[84][126],
reservoir_weight[84][127],
reservoir_weight[84][128],
reservoir_weight[84][129],
reservoir_weight[84][130],
reservoir_weight[84][131],
reservoir_weight[84][132],
reservoir_weight[84][133],
reservoir_weight[84][134],
reservoir_weight[84][135],
reservoir_weight[84][136],
reservoir_weight[84][137],
reservoir_weight[84][138],
reservoir_weight[84][139],
reservoir_weight[84][140],
reservoir_weight[84][141],
reservoir_weight[84][142],
reservoir_weight[84][143],
reservoir_weight[84][144],
reservoir_weight[84][145],
reservoir_weight[84][146],
reservoir_weight[84][147],
reservoir_weight[84][148],
reservoir_weight[84][149],
reservoir_weight[84][150],
reservoir_weight[84][151],
reservoir_weight[84][152],
reservoir_weight[84][153],
reservoir_weight[84][154],
reservoir_weight[84][155],
reservoir_weight[84][156],
reservoir_weight[84][157],
reservoir_weight[84][158],
reservoir_weight[84][159],
reservoir_weight[84][160],
reservoir_weight[84][161],
reservoir_weight[84][162],
reservoir_weight[84][163],
reservoir_weight[84][164],
reservoir_weight[84][165],
reservoir_weight[84][166],
reservoir_weight[84][167],
reservoir_weight[84][168],
reservoir_weight[84][169],
reservoir_weight[84][170],
reservoir_weight[84][171],
reservoir_weight[84][172],
reservoir_weight[84][173],
reservoir_weight[84][174],
reservoir_weight[84][175],
reservoir_weight[84][176],
reservoir_weight[84][177],
reservoir_weight[84][178],
reservoir_weight[84][179],
reservoir_weight[84][180],
reservoir_weight[84][181],
reservoir_weight[84][182],
reservoir_weight[84][183],
reservoir_weight[84][184],
reservoir_weight[84][185],
reservoir_weight[84][186],
reservoir_weight[84][187],
reservoir_weight[84][188],
reservoir_weight[84][189],
reservoir_weight[84][190],
reservoir_weight[84][191],
reservoir_weight[84][192],
reservoir_weight[84][193],
reservoir_weight[84][194],
reservoir_weight[84][195],
reservoir_weight[84][196],
reservoir_weight[84][197],
reservoir_weight[84][198],
reservoir_weight[84][199]
},
{reservoir_weight[85][0],
reservoir_weight[85][1],
reservoir_weight[85][2],
reservoir_weight[85][3],
reservoir_weight[85][4],
reservoir_weight[85][5],
reservoir_weight[85][6],
reservoir_weight[85][7],
reservoir_weight[85][8],
reservoir_weight[85][9],
reservoir_weight[85][10],
reservoir_weight[85][11],
reservoir_weight[85][12],
reservoir_weight[85][13],
reservoir_weight[85][14],
reservoir_weight[85][15],
reservoir_weight[85][16],
reservoir_weight[85][17],
reservoir_weight[85][18],
reservoir_weight[85][19],
reservoir_weight[85][20],
reservoir_weight[85][21],
reservoir_weight[85][22],
reservoir_weight[85][23],
reservoir_weight[85][24],
reservoir_weight[85][25],
reservoir_weight[85][26],
reservoir_weight[85][27],
reservoir_weight[85][28],
reservoir_weight[85][29],
reservoir_weight[85][30],
reservoir_weight[85][31],
reservoir_weight[85][32],
reservoir_weight[85][33],
reservoir_weight[85][34],
reservoir_weight[85][35],
reservoir_weight[85][36],
reservoir_weight[85][37],
reservoir_weight[85][38],
reservoir_weight[85][39],
reservoir_weight[85][40],
reservoir_weight[85][41],
reservoir_weight[85][42],
reservoir_weight[85][43],
reservoir_weight[85][44],
reservoir_weight[85][45],
reservoir_weight[85][46],
reservoir_weight[85][47],
reservoir_weight[85][48],
reservoir_weight[85][49],
reservoir_weight[85][50],
reservoir_weight[85][51],
reservoir_weight[85][52],
reservoir_weight[85][53],
reservoir_weight[85][54],
reservoir_weight[85][55],
reservoir_weight[85][56],
reservoir_weight[85][57],
reservoir_weight[85][58],
reservoir_weight[85][59],
reservoir_weight[85][60],
reservoir_weight[85][61],
reservoir_weight[85][62],
reservoir_weight[85][63],
reservoir_weight[85][64],
reservoir_weight[85][65],
reservoir_weight[85][66],
reservoir_weight[85][67],
reservoir_weight[85][68],
reservoir_weight[85][69],
reservoir_weight[85][70],
reservoir_weight[85][71],
reservoir_weight[85][72],
reservoir_weight[85][73],
reservoir_weight[85][74],
reservoir_weight[85][75],
reservoir_weight[85][76],
reservoir_weight[85][77],
reservoir_weight[85][78],
reservoir_weight[85][79],
reservoir_weight[85][80],
reservoir_weight[85][81],
reservoir_weight[85][82],
reservoir_weight[85][83],
reservoir_weight[85][84],
reservoir_weight[85][85],
reservoir_weight[85][86],
reservoir_weight[85][87],
reservoir_weight[85][88],
reservoir_weight[85][89],
reservoir_weight[85][90],
reservoir_weight[85][91],
reservoir_weight[85][92],
reservoir_weight[85][93],
reservoir_weight[85][94],
reservoir_weight[85][95],
reservoir_weight[85][96],
reservoir_weight[85][97],
reservoir_weight[85][98],
reservoir_weight[85][99],
reservoir_weight[85][100],
reservoir_weight[85][101],
reservoir_weight[85][102],
reservoir_weight[85][103],
reservoir_weight[85][104],
reservoir_weight[85][105],
reservoir_weight[85][106],
reservoir_weight[85][107],
reservoir_weight[85][108],
reservoir_weight[85][109],
reservoir_weight[85][110],
reservoir_weight[85][111],
reservoir_weight[85][112],
reservoir_weight[85][113],
reservoir_weight[85][114],
reservoir_weight[85][115],
reservoir_weight[85][116],
reservoir_weight[85][117],
reservoir_weight[85][118],
reservoir_weight[85][119],
reservoir_weight[85][120],
reservoir_weight[85][121],
reservoir_weight[85][122],
reservoir_weight[85][123],
reservoir_weight[85][124],
reservoir_weight[85][125],
reservoir_weight[85][126],
reservoir_weight[85][127],
reservoir_weight[85][128],
reservoir_weight[85][129],
reservoir_weight[85][130],
reservoir_weight[85][131],
reservoir_weight[85][132],
reservoir_weight[85][133],
reservoir_weight[85][134],
reservoir_weight[85][135],
reservoir_weight[85][136],
reservoir_weight[85][137],
reservoir_weight[85][138],
reservoir_weight[85][139],
reservoir_weight[85][140],
reservoir_weight[85][141],
reservoir_weight[85][142],
reservoir_weight[85][143],
reservoir_weight[85][144],
reservoir_weight[85][145],
reservoir_weight[85][146],
reservoir_weight[85][147],
reservoir_weight[85][148],
reservoir_weight[85][149],
reservoir_weight[85][150],
reservoir_weight[85][151],
reservoir_weight[85][152],
reservoir_weight[85][153],
reservoir_weight[85][154],
reservoir_weight[85][155],
reservoir_weight[85][156],
reservoir_weight[85][157],
reservoir_weight[85][158],
reservoir_weight[85][159],
reservoir_weight[85][160],
reservoir_weight[85][161],
reservoir_weight[85][162],
reservoir_weight[85][163],
reservoir_weight[85][164],
reservoir_weight[85][165],
reservoir_weight[85][166],
reservoir_weight[85][167],
reservoir_weight[85][168],
reservoir_weight[85][169],
reservoir_weight[85][170],
reservoir_weight[85][171],
reservoir_weight[85][172],
reservoir_weight[85][173],
reservoir_weight[85][174],
reservoir_weight[85][175],
reservoir_weight[85][176],
reservoir_weight[85][177],
reservoir_weight[85][178],
reservoir_weight[85][179],
reservoir_weight[85][180],
reservoir_weight[85][181],
reservoir_weight[85][182],
reservoir_weight[85][183],
reservoir_weight[85][184],
reservoir_weight[85][185],
reservoir_weight[85][186],
reservoir_weight[85][187],
reservoir_weight[85][188],
reservoir_weight[85][189],
reservoir_weight[85][190],
reservoir_weight[85][191],
reservoir_weight[85][192],
reservoir_weight[85][193],
reservoir_weight[85][194],
reservoir_weight[85][195],
reservoir_weight[85][196],
reservoir_weight[85][197],
reservoir_weight[85][198],
reservoir_weight[85][199]
},
{reservoir_weight[86][0],
reservoir_weight[86][1],
reservoir_weight[86][2],
reservoir_weight[86][3],
reservoir_weight[86][4],
reservoir_weight[86][5],
reservoir_weight[86][6],
reservoir_weight[86][7],
reservoir_weight[86][8],
reservoir_weight[86][9],
reservoir_weight[86][10],
reservoir_weight[86][11],
reservoir_weight[86][12],
reservoir_weight[86][13],
reservoir_weight[86][14],
reservoir_weight[86][15],
reservoir_weight[86][16],
reservoir_weight[86][17],
reservoir_weight[86][18],
reservoir_weight[86][19],
reservoir_weight[86][20],
reservoir_weight[86][21],
reservoir_weight[86][22],
reservoir_weight[86][23],
reservoir_weight[86][24],
reservoir_weight[86][25],
reservoir_weight[86][26],
reservoir_weight[86][27],
reservoir_weight[86][28],
reservoir_weight[86][29],
reservoir_weight[86][30],
reservoir_weight[86][31],
reservoir_weight[86][32],
reservoir_weight[86][33],
reservoir_weight[86][34],
reservoir_weight[86][35],
reservoir_weight[86][36],
reservoir_weight[86][37],
reservoir_weight[86][38],
reservoir_weight[86][39],
reservoir_weight[86][40],
reservoir_weight[86][41],
reservoir_weight[86][42],
reservoir_weight[86][43],
reservoir_weight[86][44],
reservoir_weight[86][45],
reservoir_weight[86][46],
reservoir_weight[86][47],
reservoir_weight[86][48],
reservoir_weight[86][49],
reservoir_weight[86][50],
reservoir_weight[86][51],
reservoir_weight[86][52],
reservoir_weight[86][53],
reservoir_weight[86][54],
reservoir_weight[86][55],
reservoir_weight[86][56],
reservoir_weight[86][57],
reservoir_weight[86][58],
reservoir_weight[86][59],
reservoir_weight[86][60],
reservoir_weight[86][61],
reservoir_weight[86][62],
reservoir_weight[86][63],
reservoir_weight[86][64],
reservoir_weight[86][65],
reservoir_weight[86][66],
reservoir_weight[86][67],
reservoir_weight[86][68],
reservoir_weight[86][69],
reservoir_weight[86][70],
reservoir_weight[86][71],
reservoir_weight[86][72],
reservoir_weight[86][73],
reservoir_weight[86][74],
reservoir_weight[86][75],
reservoir_weight[86][76],
reservoir_weight[86][77],
reservoir_weight[86][78],
reservoir_weight[86][79],
reservoir_weight[86][80],
reservoir_weight[86][81],
reservoir_weight[86][82],
reservoir_weight[86][83],
reservoir_weight[86][84],
reservoir_weight[86][85],
reservoir_weight[86][86],
reservoir_weight[86][87],
reservoir_weight[86][88],
reservoir_weight[86][89],
reservoir_weight[86][90],
reservoir_weight[86][91],
reservoir_weight[86][92],
reservoir_weight[86][93],
reservoir_weight[86][94],
reservoir_weight[86][95],
reservoir_weight[86][96],
reservoir_weight[86][97],
reservoir_weight[86][98],
reservoir_weight[86][99],
reservoir_weight[86][100],
reservoir_weight[86][101],
reservoir_weight[86][102],
reservoir_weight[86][103],
reservoir_weight[86][104],
reservoir_weight[86][105],
reservoir_weight[86][106],
reservoir_weight[86][107],
reservoir_weight[86][108],
reservoir_weight[86][109],
reservoir_weight[86][110],
reservoir_weight[86][111],
reservoir_weight[86][112],
reservoir_weight[86][113],
reservoir_weight[86][114],
reservoir_weight[86][115],
reservoir_weight[86][116],
reservoir_weight[86][117],
reservoir_weight[86][118],
reservoir_weight[86][119],
reservoir_weight[86][120],
reservoir_weight[86][121],
reservoir_weight[86][122],
reservoir_weight[86][123],
reservoir_weight[86][124],
reservoir_weight[86][125],
reservoir_weight[86][126],
reservoir_weight[86][127],
reservoir_weight[86][128],
reservoir_weight[86][129],
reservoir_weight[86][130],
reservoir_weight[86][131],
reservoir_weight[86][132],
reservoir_weight[86][133],
reservoir_weight[86][134],
reservoir_weight[86][135],
reservoir_weight[86][136],
reservoir_weight[86][137],
reservoir_weight[86][138],
reservoir_weight[86][139],
reservoir_weight[86][140],
reservoir_weight[86][141],
reservoir_weight[86][142],
reservoir_weight[86][143],
reservoir_weight[86][144],
reservoir_weight[86][145],
reservoir_weight[86][146],
reservoir_weight[86][147],
reservoir_weight[86][148],
reservoir_weight[86][149],
reservoir_weight[86][150],
reservoir_weight[86][151],
reservoir_weight[86][152],
reservoir_weight[86][153],
reservoir_weight[86][154],
reservoir_weight[86][155],
reservoir_weight[86][156],
reservoir_weight[86][157],
reservoir_weight[86][158],
reservoir_weight[86][159],
reservoir_weight[86][160],
reservoir_weight[86][161],
reservoir_weight[86][162],
reservoir_weight[86][163],
reservoir_weight[86][164],
reservoir_weight[86][165],
reservoir_weight[86][166],
reservoir_weight[86][167],
reservoir_weight[86][168],
reservoir_weight[86][169],
reservoir_weight[86][170],
reservoir_weight[86][171],
reservoir_weight[86][172],
reservoir_weight[86][173],
reservoir_weight[86][174],
reservoir_weight[86][175],
reservoir_weight[86][176],
reservoir_weight[86][177],
reservoir_weight[86][178],
reservoir_weight[86][179],
reservoir_weight[86][180],
reservoir_weight[86][181],
reservoir_weight[86][182],
reservoir_weight[86][183],
reservoir_weight[86][184],
reservoir_weight[86][185],
reservoir_weight[86][186],
reservoir_weight[86][187],
reservoir_weight[86][188],
reservoir_weight[86][189],
reservoir_weight[86][190],
reservoir_weight[86][191],
reservoir_weight[86][192],
reservoir_weight[86][193],
reservoir_weight[86][194],
reservoir_weight[86][195],
reservoir_weight[86][196],
reservoir_weight[86][197],
reservoir_weight[86][198],
reservoir_weight[86][199]
},
{reservoir_weight[87][0],
reservoir_weight[87][1],
reservoir_weight[87][2],
reservoir_weight[87][3],
reservoir_weight[87][4],
reservoir_weight[87][5],
reservoir_weight[87][6],
reservoir_weight[87][7],
reservoir_weight[87][8],
reservoir_weight[87][9],
reservoir_weight[87][10],
reservoir_weight[87][11],
reservoir_weight[87][12],
reservoir_weight[87][13],
reservoir_weight[87][14],
reservoir_weight[87][15],
reservoir_weight[87][16],
reservoir_weight[87][17],
reservoir_weight[87][18],
reservoir_weight[87][19],
reservoir_weight[87][20],
reservoir_weight[87][21],
reservoir_weight[87][22],
reservoir_weight[87][23],
reservoir_weight[87][24],
reservoir_weight[87][25],
reservoir_weight[87][26],
reservoir_weight[87][27],
reservoir_weight[87][28],
reservoir_weight[87][29],
reservoir_weight[87][30],
reservoir_weight[87][31],
reservoir_weight[87][32],
reservoir_weight[87][33],
reservoir_weight[87][34],
reservoir_weight[87][35],
reservoir_weight[87][36],
reservoir_weight[87][37],
reservoir_weight[87][38],
reservoir_weight[87][39],
reservoir_weight[87][40],
reservoir_weight[87][41],
reservoir_weight[87][42],
reservoir_weight[87][43],
reservoir_weight[87][44],
reservoir_weight[87][45],
reservoir_weight[87][46],
reservoir_weight[87][47],
reservoir_weight[87][48],
reservoir_weight[87][49],
reservoir_weight[87][50],
reservoir_weight[87][51],
reservoir_weight[87][52],
reservoir_weight[87][53],
reservoir_weight[87][54],
reservoir_weight[87][55],
reservoir_weight[87][56],
reservoir_weight[87][57],
reservoir_weight[87][58],
reservoir_weight[87][59],
reservoir_weight[87][60],
reservoir_weight[87][61],
reservoir_weight[87][62],
reservoir_weight[87][63],
reservoir_weight[87][64],
reservoir_weight[87][65],
reservoir_weight[87][66],
reservoir_weight[87][67],
reservoir_weight[87][68],
reservoir_weight[87][69],
reservoir_weight[87][70],
reservoir_weight[87][71],
reservoir_weight[87][72],
reservoir_weight[87][73],
reservoir_weight[87][74],
reservoir_weight[87][75],
reservoir_weight[87][76],
reservoir_weight[87][77],
reservoir_weight[87][78],
reservoir_weight[87][79],
reservoir_weight[87][80],
reservoir_weight[87][81],
reservoir_weight[87][82],
reservoir_weight[87][83],
reservoir_weight[87][84],
reservoir_weight[87][85],
reservoir_weight[87][86],
reservoir_weight[87][87],
reservoir_weight[87][88],
reservoir_weight[87][89],
reservoir_weight[87][90],
reservoir_weight[87][91],
reservoir_weight[87][92],
reservoir_weight[87][93],
reservoir_weight[87][94],
reservoir_weight[87][95],
reservoir_weight[87][96],
reservoir_weight[87][97],
reservoir_weight[87][98],
reservoir_weight[87][99],
reservoir_weight[87][100],
reservoir_weight[87][101],
reservoir_weight[87][102],
reservoir_weight[87][103],
reservoir_weight[87][104],
reservoir_weight[87][105],
reservoir_weight[87][106],
reservoir_weight[87][107],
reservoir_weight[87][108],
reservoir_weight[87][109],
reservoir_weight[87][110],
reservoir_weight[87][111],
reservoir_weight[87][112],
reservoir_weight[87][113],
reservoir_weight[87][114],
reservoir_weight[87][115],
reservoir_weight[87][116],
reservoir_weight[87][117],
reservoir_weight[87][118],
reservoir_weight[87][119],
reservoir_weight[87][120],
reservoir_weight[87][121],
reservoir_weight[87][122],
reservoir_weight[87][123],
reservoir_weight[87][124],
reservoir_weight[87][125],
reservoir_weight[87][126],
reservoir_weight[87][127],
reservoir_weight[87][128],
reservoir_weight[87][129],
reservoir_weight[87][130],
reservoir_weight[87][131],
reservoir_weight[87][132],
reservoir_weight[87][133],
reservoir_weight[87][134],
reservoir_weight[87][135],
reservoir_weight[87][136],
reservoir_weight[87][137],
reservoir_weight[87][138],
reservoir_weight[87][139],
reservoir_weight[87][140],
reservoir_weight[87][141],
reservoir_weight[87][142],
reservoir_weight[87][143],
reservoir_weight[87][144],
reservoir_weight[87][145],
reservoir_weight[87][146],
reservoir_weight[87][147],
reservoir_weight[87][148],
reservoir_weight[87][149],
reservoir_weight[87][150],
reservoir_weight[87][151],
reservoir_weight[87][152],
reservoir_weight[87][153],
reservoir_weight[87][154],
reservoir_weight[87][155],
reservoir_weight[87][156],
reservoir_weight[87][157],
reservoir_weight[87][158],
reservoir_weight[87][159],
reservoir_weight[87][160],
reservoir_weight[87][161],
reservoir_weight[87][162],
reservoir_weight[87][163],
reservoir_weight[87][164],
reservoir_weight[87][165],
reservoir_weight[87][166],
reservoir_weight[87][167],
reservoir_weight[87][168],
reservoir_weight[87][169],
reservoir_weight[87][170],
reservoir_weight[87][171],
reservoir_weight[87][172],
reservoir_weight[87][173],
reservoir_weight[87][174],
reservoir_weight[87][175],
reservoir_weight[87][176],
reservoir_weight[87][177],
reservoir_weight[87][178],
reservoir_weight[87][179],
reservoir_weight[87][180],
reservoir_weight[87][181],
reservoir_weight[87][182],
reservoir_weight[87][183],
reservoir_weight[87][184],
reservoir_weight[87][185],
reservoir_weight[87][186],
reservoir_weight[87][187],
reservoir_weight[87][188],
reservoir_weight[87][189],
reservoir_weight[87][190],
reservoir_weight[87][191],
reservoir_weight[87][192],
reservoir_weight[87][193],
reservoir_weight[87][194],
reservoir_weight[87][195],
reservoir_weight[87][196],
reservoir_weight[87][197],
reservoir_weight[87][198],
reservoir_weight[87][199]
},
{reservoir_weight[88][0],
reservoir_weight[88][1],
reservoir_weight[88][2],
reservoir_weight[88][3],
reservoir_weight[88][4],
reservoir_weight[88][5],
reservoir_weight[88][6],
reservoir_weight[88][7],
reservoir_weight[88][8],
reservoir_weight[88][9],
reservoir_weight[88][10],
reservoir_weight[88][11],
reservoir_weight[88][12],
reservoir_weight[88][13],
reservoir_weight[88][14],
reservoir_weight[88][15],
reservoir_weight[88][16],
reservoir_weight[88][17],
reservoir_weight[88][18],
reservoir_weight[88][19],
reservoir_weight[88][20],
reservoir_weight[88][21],
reservoir_weight[88][22],
reservoir_weight[88][23],
reservoir_weight[88][24],
reservoir_weight[88][25],
reservoir_weight[88][26],
reservoir_weight[88][27],
reservoir_weight[88][28],
reservoir_weight[88][29],
reservoir_weight[88][30],
reservoir_weight[88][31],
reservoir_weight[88][32],
reservoir_weight[88][33],
reservoir_weight[88][34],
reservoir_weight[88][35],
reservoir_weight[88][36],
reservoir_weight[88][37],
reservoir_weight[88][38],
reservoir_weight[88][39],
reservoir_weight[88][40],
reservoir_weight[88][41],
reservoir_weight[88][42],
reservoir_weight[88][43],
reservoir_weight[88][44],
reservoir_weight[88][45],
reservoir_weight[88][46],
reservoir_weight[88][47],
reservoir_weight[88][48],
reservoir_weight[88][49],
reservoir_weight[88][50],
reservoir_weight[88][51],
reservoir_weight[88][52],
reservoir_weight[88][53],
reservoir_weight[88][54],
reservoir_weight[88][55],
reservoir_weight[88][56],
reservoir_weight[88][57],
reservoir_weight[88][58],
reservoir_weight[88][59],
reservoir_weight[88][60],
reservoir_weight[88][61],
reservoir_weight[88][62],
reservoir_weight[88][63],
reservoir_weight[88][64],
reservoir_weight[88][65],
reservoir_weight[88][66],
reservoir_weight[88][67],
reservoir_weight[88][68],
reservoir_weight[88][69],
reservoir_weight[88][70],
reservoir_weight[88][71],
reservoir_weight[88][72],
reservoir_weight[88][73],
reservoir_weight[88][74],
reservoir_weight[88][75],
reservoir_weight[88][76],
reservoir_weight[88][77],
reservoir_weight[88][78],
reservoir_weight[88][79],
reservoir_weight[88][80],
reservoir_weight[88][81],
reservoir_weight[88][82],
reservoir_weight[88][83],
reservoir_weight[88][84],
reservoir_weight[88][85],
reservoir_weight[88][86],
reservoir_weight[88][87],
reservoir_weight[88][88],
reservoir_weight[88][89],
reservoir_weight[88][90],
reservoir_weight[88][91],
reservoir_weight[88][92],
reservoir_weight[88][93],
reservoir_weight[88][94],
reservoir_weight[88][95],
reservoir_weight[88][96],
reservoir_weight[88][97],
reservoir_weight[88][98],
reservoir_weight[88][99],
reservoir_weight[88][100],
reservoir_weight[88][101],
reservoir_weight[88][102],
reservoir_weight[88][103],
reservoir_weight[88][104],
reservoir_weight[88][105],
reservoir_weight[88][106],
reservoir_weight[88][107],
reservoir_weight[88][108],
reservoir_weight[88][109],
reservoir_weight[88][110],
reservoir_weight[88][111],
reservoir_weight[88][112],
reservoir_weight[88][113],
reservoir_weight[88][114],
reservoir_weight[88][115],
reservoir_weight[88][116],
reservoir_weight[88][117],
reservoir_weight[88][118],
reservoir_weight[88][119],
reservoir_weight[88][120],
reservoir_weight[88][121],
reservoir_weight[88][122],
reservoir_weight[88][123],
reservoir_weight[88][124],
reservoir_weight[88][125],
reservoir_weight[88][126],
reservoir_weight[88][127],
reservoir_weight[88][128],
reservoir_weight[88][129],
reservoir_weight[88][130],
reservoir_weight[88][131],
reservoir_weight[88][132],
reservoir_weight[88][133],
reservoir_weight[88][134],
reservoir_weight[88][135],
reservoir_weight[88][136],
reservoir_weight[88][137],
reservoir_weight[88][138],
reservoir_weight[88][139],
reservoir_weight[88][140],
reservoir_weight[88][141],
reservoir_weight[88][142],
reservoir_weight[88][143],
reservoir_weight[88][144],
reservoir_weight[88][145],
reservoir_weight[88][146],
reservoir_weight[88][147],
reservoir_weight[88][148],
reservoir_weight[88][149],
reservoir_weight[88][150],
reservoir_weight[88][151],
reservoir_weight[88][152],
reservoir_weight[88][153],
reservoir_weight[88][154],
reservoir_weight[88][155],
reservoir_weight[88][156],
reservoir_weight[88][157],
reservoir_weight[88][158],
reservoir_weight[88][159],
reservoir_weight[88][160],
reservoir_weight[88][161],
reservoir_weight[88][162],
reservoir_weight[88][163],
reservoir_weight[88][164],
reservoir_weight[88][165],
reservoir_weight[88][166],
reservoir_weight[88][167],
reservoir_weight[88][168],
reservoir_weight[88][169],
reservoir_weight[88][170],
reservoir_weight[88][171],
reservoir_weight[88][172],
reservoir_weight[88][173],
reservoir_weight[88][174],
reservoir_weight[88][175],
reservoir_weight[88][176],
reservoir_weight[88][177],
reservoir_weight[88][178],
reservoir_weight[88][179],
reservoir_weight[88][180],
reservoir_weight[88][181],
reservoir_weight[88][182],
reservoir_weight[88][183],
reservoir_weight[88][184],
reservoir_weight[88][185],
reservoir_weight[88][186],
reservoir_weight[88][187],
reservoir_weight[88][188],
reservoir_weight[88][189],
reservoir_weight[88][190],
reservoir_weight[88][191],
reservoir_weight[88][192],
reservoir_weight[88][193],
reservoir_weight[88][194],
reservoir_weight[88][195],
reservoir_weight[88][196],
reservoir_weight[88][197],
reservoir_weight[88][198],
reservoir_weight[88][199]
},
{reservoir_weight[89][0],
reservoir_weight[89][1],
reservoir_weight[89][2],
reservoir_weight[89][3],
reservoir_weight[89][4],
reservoir_weight[89][5],
reservoir_weight[89][6],
reservoir_weight[89][7],
reservoir_weight[89][8],
reservoir_weight[89][9],
reservoir_weight[89][10],
reservoir_weight[89][11],
reservoir_weight[89][12],
reservoir_weight[89][13],
reservoir_weight[89][14],
reservoir_weight[89][15],
reservoir_weight[89][16],
reservoir_weight[89][17],
reservoir_weight[89][18],
reservoir_weight[89][19],
reservoir_weight[89][20],
reservoir_weight[89][21],
reservoir_weight[89][22],
reservoir_weight[89][23],
reservoir_weight[89][24],
reservoir_weight[89][25],
reservoir_weight[89][26],
reservoir_weight[89][27],
reservoir_weight[89][28],
reservoir_weight[89][29],
reservoir_weight[89][30],
reservoir_weight[89][31],
reservoir_weight[89][32],
reservoir_weight[89][33],
reservoir_weight[89][34],
reservoir_weight[89][35],
reservoir_weight[89][36],
reservoir_weight[89][37],
reservoir_weight[89][38],
reservoir_weight[89][39],
reservoir_weight[89][40],
reservoir_weight[89][41],
reservoir_weight[89][42],
reservoir_weight[89][43],
reservoir_weight[89][44],
reservoir_weight[89][45],
reservoir_weight[89][46],
reservoir_weight[89][47],
reservoir_weight[89][48],
reservoir_weight[89][49],
reservoir_weight[89][50],
reservoir_weight[89][51],
reservoir_weight[89][52],
reservoir_weight[89][53],
reservoir_weight[89][54],
reservoir_weight[89][55],
reservoir_weight[89][56],
reservoir_weight[89][57],
reservoir_weight[89][58],
reservoir_weight[89][59],
reservoir_weight[89][60],
reservoir_weight[89][61],
reservoir_weight[89][62],
reservoir_weight[89][63],
reservoir_weight[89][64],
reservoir_weight[89][65],
reservoir_weight[89][66],
reservoir_weight[89][67],
reservoir_weight[89][68],
reservoir_weight[89][69],
reservoir_weight[89][70],
reservoir_weight[89][71],
reservoir_weight[89][72],
reservoir_weight[89][73],
reservoir_weight[89][74],
reservoir_weight[89][75],
reservoir_weight[89][76],
reservoir_weight[89][77],
reservoir_weight[89][78],
reservoir_weight[89][79],
reservoir_weight[89][80],
reservoir_weight[89][81],
reservoir_weight[89][82],
reservoir_weight[89][83],
reservoir_weight[89][84],
reservoir_weight[89][85],
reservoir_weight[89][86],
reservoir_weight[89][87],
reservoir_weight[89][88],
reservoir_weight[89][89],
reservoir_weight[89][90],
reservoir_weight[89][91],
reservoir_weight[89][92],
reservoir_weight[89][93],
reservoir_weight[89][94],
reservoir_weight[89][95],
reservoir_weight[89][96],
reservoir_weight[89][97],
reservoir_weight[89][98],
reservoir_weight[89][99],
reservoir_weight[89][100],
reservoir_weight[89][101],
reservoir_weight[89][102],
reservoir_weight[89][103],
reservoir_weight[89][104],
reservoir_weight[89][105],
reservoir_weight[89][106],
reservoir_weight[89][107],
reservoir_weight[89][108],
reservoir_weight[89][109],
reservoir_weight[89][110],
reservoir_weight[89][111],
reservoir_weight[89][112],
reservoir_weight[89][113],
reservoir_weight[89][114],
reservoir_weight[89][115],
reservoir_weight[89][116],
reservoir_weight[89][117],
reservoir_weight[89][118],
reservoir_weight[89][119],
reservoir_weight[89][120],
reservoir_weight[89][121],
reservoir_weight[89][122],
reservoir_weight[89][123],
reservoir_weight[89][124],
reservoir_weight[89][125],
reservoir_weight[89][126],
reservoir_weight[89][127],
reservoir_weight[89][128],
reservoir_weight[89][129],
reservoir_weight[89][130],
reservoir_weight[89][131],
reservoir_weight[89][132],
reservoir_weight[89][133],
reservoir_weight[89][134],
reservoir_weight[89][135],
reservoir_weight[89][136],
reservoir_weight[89][137],
reservoir_weight[89][138],
reservoir_weight[89][139],
reservoir_weight[89][140],
reservoir_weight[89][141],
reservoir_weight[89][142],
reservoir_weight[89][143],
reservoir_weight[89][144],
reservoir_weight[89][145],
reservoir_weight[89][146],
reservoir_weight[89][147],
reservoir_weight[89][148],
reservoir_weight[89][149],
reservoir_weight[89][150],
reservoir_weight[89][151],
reservoir_weight[89][152],
reservoir_weight[89][153],
reservoir_weight[89][154],
reservoir_weight[89][155],
reservoir_weight[89][156],
reservoir_weight[89][157],
reservoir_weight[89][158],
reservoir_weight[89][159],
reservoir_weight[89][160],
reservoir_weight[89][161],
reservoir_weight[89][162],
reservoir_weight[89][163],
reservoir_weight[89][164],
reservoir_weight[89][165],
reservoir_weight[89][166],
reservoir_weight[89][167],
reservoir_weight[89][168],
reservoir_weight[89][169],
reservoir_weight[89][170],
reservoir_weight[89][171],
reservoir_weight[89][172],
reservoir_weight[89][173],
reservoir_weight[89][174],
reservoir_weight[89][175],
reservoir_weight[89][176],
reservoir_weight[89][177],
reservoir_weight[89][178],
reservoir_weight[89][179],
reservoir_weight[89][180],
reservoir_weight[89][181],
reservoir_weight[89][182],
reservoir_weight[89][183],
reservoir_weight[89][184],
reservoir_weight[89][185],
reservoir_weight[89][186],
reservoir_weight[89][187],
reservoir_weight[89][188],
reservoir_weight[89][189],
reservoir_weight[89][190],
reservoir_weight[89][191],
reservoir_weight[89][192],
reservoir_weight[89][193],
reservoir_weight[89][194],
reservoir_weight[89][195],
reservoir_weight[89][196],
reservoir_weight[89][197],
reservoir_weight[89][198],
reservoir_weight[89][199]
},
{reservoir_weight[90][0],
reservoir_weight[90][1],
reservoir_weight[90][2],
reservoir_weight[90][3],
reservoir_weight[90][4],
reservoir_weight[90][5],
reservoir_weight[90][6],
reservoir_weight[90][7],
reservoir_weight[90][8],
reservoir_weight[90][9],
reservoir_weight[90][10],
reservoir_weight[90][11],
reservoir_weight[90][12],
reservoir_weight[90][13],
reservoir_weight[90][14],
reservoir_weight[90][15],
reservoir_weight[90][16],
reservoir_weight[90][17],
reservoir_weight[90][18],
reservoir_weight[90][19],
reservoir_weight[90][20],
reservoir_weight[90][21],
reservoir_weight[90][22],
reservoir_weight[90][23],
reservoir_weight[90][24],
reservoir_weight[90][25],
reservoir_weight[90][26],
reservoir_weight[90][27],
reservoir_weight[90][28],
reservoir_weight[90][29],
reservoir_weight[90][30],
reservoir_weight[90][31],
reservoir_weight[90][32],
reservoir_weight[90][33],
reservoir_weight[90][34],
reservoir_weight[90][35],
reservoir_weight[90][36],
reservoir_weight[90][37],
reservoir_weight[90][38],
reservoir_weight[90][39],
reservoir_weight[90][40],
reservoir_weight[90][41],
reservoir_weight[90][42],
reservoir_weight[90][43],
reservoir_weight[90][44],
reservoir_weight[90][45],
reservoir_weight[90][46],
reservoir_weight[90][47],
reservoir_weight[90][48],
reservoir_weight[90][49],
reservoir_weight[90][50],
reservoir_weight[90][51],
reservoir_weight[90][52],
reservoir_weight[90][53],
reservoir_weight[90][54],
reservoir_weight[90][55],
reservoir_weight[90][56],
reservoir_weight[90][57],
reservoir_weight[90][58],
reservoir_weight[90][59],
reservoir_weight[90][60],
reservoir_weight[90][61],
reservoir_weight[90][62],
reservoir_weight[90][63],
reservoir_weight[90][64],
reservoir_weight[90][65],
reservoir_weight[90][66],
reservoir_weight[90][67],
reservoir_weight[90][68],
reservoir_weight[90][69],
reservoir_weight[90][70],
reservoir_weight[90][71],
reservoir_weight[90][72],
reservoir_weight[90][73],
reservoir_weight[90][74],
reservoir_weight[90][75],
reservoir_weight[90][76],
reservoir_weight[90][77],
reservoir_weight[90][78],
reservoir_weight[90][79],
reservoir_weight[90][80],
reservoir_weight[90][81],
reservoir_weight[90][82],
reservoir_weight[90][83],
reservoir_weight[90][84],
reservoir_weight[90][85],
reservoir_weight[90][86],
reservoir_weight[90][87],
reservoir_weight[90][88],
reservoir_weight[90][89],
reservoir_weight[90][90],
reservoir_weight[90][91],
reservoir_weight[90][92],
reservoir_weight[90][93],
reservoir_weight[90][94],
reservoir_weight[90][95],
reservoir_weight[90][96],
reservoir_weight[90][97],
reservoir_weight[90][98],
reservoir_weight[90][99],
reservoir_weight[90][100],
reservoir_weight[90][101],
reservoir_weight[90][102],
reservoir_weight[90][103],
reservoir_weight[90][104],
reservoir_weight[90][105],
reservoir_weight[90][106],
reservoir_weight[90][107],
reservoir_weight[90][108],
reservoir_weight[90][109],
reservoir_weight[90][110],
reservoir_weight[90][111],
reservoir_weight[90][112],
reservoir_weight[90][113],
reservoir_weight[90][114],
reservoir_weight[90][115],
reservoir_weight[90][116],
reservoir_weight[90][117],
reservoir_weight[90][118],
reservoir_weight[90][119],
reservoir_weight[90][120],
reservoir_weight[90][121],
reservoir_weight[90][122],
reservoir_weight[90][123],
reservoir_weight[90][124],
reservoir_weight[90][125],
reservoir_weight[90][126],
reservoir_weight[90][127],
reservoir_weight[90][128],
reservoir_weight[90][129],
reservoir_weight[90][130],
reservoir_weight[90][131],
reservoir_weight[90][132],
reservoir_weight[90][133],
reservoir_weight[90][134],
reservoir_weight[90][135],
reservoir_weight[90][136],
reservoir_weight[90][137],
reservoir_weight[90][138],
reservoir_weight[90][139],
reservoir_weight[90][140],
reservoir_weight[90][141],
reservoir_weight[90][142],
reservoir_weight[90][143],
reservoir_weight[90][144],
reservoir_weight[90][145],
reservoir_weight[90][146],
reservoir_weight[90][147],
reservoir_weight[90][148],
reservoir_weight[90][149],
reservoir_weight[90][150],
reservoir_weight[90][151],
reservoir_weight[90][152],
reservoir_weight[90][153],
reservoir_weight[90][154],
reservoir_weight[90][155],
reservoir_weight[90][156],
reservoir_weight[90][157],
reservoir_weight[90][158],
reservoir_weight[90][159],
reservoir_weight[90][160],
reservoir_weight[90][161],
reservoir_weight[90][162],
reservoir_weight[90][163],
reservoir_weight[90][164],
reservoir_weight[90][165],
reservoir_weight[90][166],
reservoir_weight[90][167],
reservoir_weight[90][168],
reservoir_weight[90][169],
reservoir_weight[90][170],
reservoir_weight[90][171],
reservoir_weight[90][172],
reservoir_weight[90][173],
reservoir_weight[90][174],
reservoir_weight[90][175],
reservoir_weight[90][176],
reservoir_weight[90][177],
reservoir_weight[90][178],
reservoir_weight[90][179],
reservoir_weight[90][180],
reservoir_weight[90][181],
reservoir_weight[90][182],
reservoir_weight[90][183],
reservoir_weight[90][184],
reservoir_weight[90][185],
reservoir_weight[90][186],
reservoir_weight[90][187],
reservoir_weight[90][188],
reservoir_weight[90][189],
reservoir_weight[90][190],
reservoir_weight[90][191],
reservoir_weight[90][192],
reservoir_weight[90][193],
reservoir_weight[90][194],
reservoir_weight[90][195],
reservoir_weight[90][196],
reservoir_weight[90][197],
reservoir_weight[90][198],
reservoir_weight[90][199]
},
{reservoir_weight[91][0],
reservoir_weight[91][1],
reservoir_weight[91][2],
reservoir_weight[91][3],
reservoir_weight[91][4],
reservoir_weight[91][5],
reservoir_weight[91][6],
reservoir_weight[91][7],
reservoir_weight[91][8],
reservoir_weight[91][9],
reservoir_weight[91][10],
reservoir_weight[91][11],
reservoir_weight[91][12],
reservoir_weight[91][13],
reservoir_weight[91][14],
reservoir_weight[91][15],
reservoir_weight[91][16],
reservoir_weight[91][17],
reservoir_weight[91][18],
reservoir_weight[91][19],
reservoir_weight[91][20],
reservoir_weight[91][21],
reservoir_weight[91][22],
reservoir_weight[91][23],
reservoir_weight[91][24],
reservoir_weight[91][25],
reservoir_weight[91][26],
reservoir_weight[91][27],
reservoir_weight[91][28],
reservoir_weight[91][29],
reservoir_weight[91][30],
reservoir_weight[91][31],
reservoir_weight[91][32],
reservoir_weight[91][33],
reservoir_weight[91][34],
reservoir_weight[91][35],
reservoir_weight[91][36],
reservoir_weight[91][37],
reservoir_weight[91][38],
reservoir_weight[91][39],
reservoir_weight[91][40],
reservoir_weight[91][41],
reservoir_weight[91][42],
reservoir_weight[91][43],
reservoir_weight[91][44],
reservoir_weight[91][45],
reservoir_weight[91][46],
reservoir_weight[91][47],
reservoir_weight[91][48],
reservoir_weight[91][49],
reservoir_weight[91][50],
reservoir_weight[91][51],
reservoir_weight[91][52],
reservoir_weight[91][53],
reservoir_weight[91][54],
reservoir_weight[91][55],
reservoir_weight[91][56],
reservoir_weight[91][57],
reservoir_weight[91][58],
reservoir_weight[91][59],
reservoir_weight[91][60],
reservoir_weight[91][61],
reservoir_weight[91][62],
reservoir_weight[91][63],
reservoir_weight[91][64],
reservoir_weight[91][65],
reservoir_weight[91][66],
reservoir_weight[91][67],
reservoir_weight[91][68],
reservoir_weight[91][69],
reservoir_weight[91][70],
reservoir_weight[91][71],
reservoir_weight[91][72],
reservoir_weight[91][73],
reservoir_weight[91][74],
reservoir_weight[91][75],
reservoir_weight[91][76],
reservoir_weight[91][77],
reservoir_weight[91][78],
reservoir_weight[91][79],
reservoir_weight[91][80],
reservoir_weight[91][81],
reservoir_weight[91][82],
reservoir_weight[91][83],
reservoir_weight[91][84],
reservoir_weight[91][85],
reservoir_weight[91][86],
reservoir_weight[91][87],
reservoir_weight[91][88],
reservoir_weight[91][89],
reservoir_weight[91][90],
reservoir_weight[91][91],
reservoir_weight[91][92],
reservoir_weight[91][93],
reservoir_weight[91][94],
reservoir_weight[91][95],
reservoir_weight[91][96],
reservoir_weight[91][97],
reservoir_weight[91][98],
reservoir_weight[91][99],
reservoir_weight[91][100],
reservoir_weight[91][101],
reservoir_weight[91][102],
reservoir_weight[91][103],
reservoir_weight[91][104],
reservoir_weight[91][105],
reservoir_weight[91][106],
reservoir_weight[91][107],
reservoir_weight[91][108],
reservoir_weight[91][109],
reservoir_weight[91][110],
reservoir_weight[91][111],
reservoir_weight[91][112],
reservoir_weight[91][113],
reservoir_weight[91][114],
reservoir_weight[91][115],
reservoir_weight[91][116],
reservoir_weight[91][117],
reservoir_weight[91][118],
reservoir_weight[91][119],
reservoir_weight[91][120],
reservoir_weight[91][121],
reservoir_weight[91][122],
reservoir_weight[91][123],
reservoir_weight[91][124],
reservoir_weight[91][125],
reservoir_weight[91][126],
reservoir_weight[91][127],
reservoir_weight[91][128],
reservoir_weight[91][129],
reservoir_weight[91][130],
reservoir_weight[91][131],
reservoir_weight[91][132],
reservoir_weight[91][133],
reservoir_weight[91][134],
reservoir_weight[91][135],
reservoir_weight[91][136],
reservoir_weight[91][137],
reservoir_weight[91][138],
reservoir_weight[91][139],
reservoir_weight[91][140],
reservoir_weight[91][141],
reservoir_weight[91][142],
reservoir_weight[91][143],
reservoir_weight[91][144],
reservoir_weight[91][145],
reservoir_weight[91][146],
reservoir_weight[91][147],
reservoir_weight[91][148],
reservoir_weight[91][149],
reservoir_weight[91][150],
reservoir_weight[91][151],
reservoir_weight[91][152],
reservoir_weight[91][153],
reservoir_weight[91][154],
reservoir_weight[91][155],
reservoir_weight[91][156],
reservoir_weight[91][157],
reservoir_weight[91][158],
reservoir_weight[91][159],
reservoir_weight[91][160],
reservoir_weight[91][161],
reservoir_weight[91][162],
reservoir_weight[91][163],
reservoir_weight[91][164],
reservoir_weight[91][165],
reservoir_weight[91][166],
reservoir_weight[91][167],
reservoir_weight[91][168],
reservoir_weight[91][169],
reservoir_weight[91][170],
reservoir_weight[91][171],
reservoir_weight[91][172],
reservoir_weight[91][173],
reservoir_weight[91][174],
reservoir_weight[91][175],
reservoir_weight[91][176],
reservoir_weight[91][177],
reservoir_weight[91][178],
reservoir_weight[91][179],
reservoir_weight[91][180],
reservoir_weight[91][181],
reservoir_weight[91][182],
reservoir_weight[91][183],
reservoir_weight[91][184],
reservoir_weight[91][185],
reservoir_weight[91][186],
reservoir_weight[91][187],
reservoir_weight[91][188],
reservoir_weight[91][189],
reservoir_weight[91][190],
reservoir_weight[91][191],
reservoir_weight[91][192],
reservoir_weight[91][193],
reservoir_weight[91][194],
reservoir_weight[91][195],
reservoir_weight[91][196],
reservoir_weight[91][197],
reservoir_weight[91][198],
reservoir_weight[91][199]
},
{reservoir_weight[92][0],
reservoir_weight[92][1],
reservoir_weight[92][2],
reservoir_weight[92][3],
reservoir_weight[92][4],
reservoir_weight[92][5],
reservoir_weight[92][6],
reservoir_weight[92][7],
reservoir_weight[92][8],
reservoir_weight[92][9],
reservoir_weight[92][10],
reservoir_weight[92][11],
reservoir_weight[92][12],
reservoir_weight[92][13],
reservoir_weight[92][14],
reservoir_weight[92][15],
reservoir_weight[92][16],
reservoir_weight[92][17],
reservoir_weight[92][18],
reservoir_weight[92][19],
reservoir_weight[92][20],
reservoir_weight[92][21],
reservoir_weight[92][22],
reservoir_weight[92][23],
reservoir_weight[92][24],
reservoir_weight[92][25],
reservoir_weight[92][26],
reservoir_weight[92][27],
reservoir_weight[92][28],
reservoir_weight[92][29],
reservoir_weight[92][30],
reservoir_weight[92][31],
reservoir_weight[92][32],
reservoir_weight[92][33],
reservoir_weight[92][34],
reservoir_weight[92][35],
reservoir_weight[92][36],
reservoir_weight[92][37],
reservoir_weight[92][38],
reservoir_weight[92][39],
reservoir_weight[92][40],
reservoir_weight[92][41],
reservoir_weight[92][42],
reservoir_weight[92][43],
reservoir_weight[92][44],
reservoir_weight[92][45],
reservoir_weight[92][46],
reservoir_weight[92][47],
reservoir_weight[92][48],
reservoir_weight[92][49],
reservoir_weight[92][50],
reservoir_weight[92][51],
reservoir_weight[92][52],
reservoir_weight[92][53],
reservoir_weight[92][54],
reservoir_weight[92][55],
reservoir_weight[92][56],
reservoir_weight[92][57],
reservoir_weight[92][58],
reservoir_weight[92][59],
reservoir_weight[92][60],
reservoir_weight[92][61],
reservoir_weight[92][62],
reservoir_weight[92][63],
reservoir_weight[92][64],
reservoir_weight[92][65],
reservoir_weight[92][66],
reservoir_weight[92][67],
reservoir_weight[92][68],
reservoir_weight[92][69],
reservoir_weight[92][70],
reservoir_weight[92][71],
reservoir_weight[92][72],
reservoir_weight[92][73],
reservoir_weight[92][74],
reservoir_weight[92][75],
reservoir_weight[92][76],
reservoir_weight[92][77],
reservoir_weight[92][78],
reservoir_weight[92][79],
reservoir_weight[92][80],
reservoir_weight[92][81],
reservoir_weight[92][82],
reservoir_weight[92][83],
reservoir_weight[92][84],
reservoir_weight[92][85],
reservoir_weight[92][86],
reservoir_weight[92][87],
reservoir_weight[92][88],
reservoir_weight[92][89],
reservoir_weight[92][90],
reservoir_weight[92][91],
reservoir_weight[92][92],
reservoir_weight[92][93],
reservoir_weight[92][94],
reservoir_weight[92][95],
reservoir_weight[92][96],
reservoir_weight[92][97],
reservoir_weight[92][98],
reservoir_weight[92][99],
reservoir_weight[92][100],
reservoir_weight[92][101],
reservoir_weight[92][102],
reservoir_weight[92][103],
reservoir_weight[92][104],
reservoir_weight[92][105],
reservoir_weight[92][106],
reservoir_weight[92][107],
reservoir_weight[92][108],
reservoir_weight[92][109],
reservoir_weight[92][110],
reservoir_weight[92][111],
reservoir_weight[92][112],
reservoir_weight[92][113],
reservoir_weight[92][114],
reservoir_weight[92][115],
reservoir_weight[92][116],
reservoir_weight[92][117],
reservoir_weight[92][118],
reservoir_weight[92][119],
reservoir_weight[92][120],
reservoir_weight[92][121],
reservoir_weight[92][122],
reservoir_weight[92][123],
reservoir_weight[92][124],
reservoir_weight[92][125],
reservoir_weight[92][126],
reservoir_weight[92][127],
reservoir_weight[92][128],
reservoir_weight[92][129],
reservoir_weight[92][130],
reservoir_weight[92][131],
reservoir_weight[92][132],
reservoir_weight[92][133],
reservoir_weight[92][134],
reservoir_weight[92][135],
reservoir_weight[92][136],
reservoir_weight[92][137],
reservoir_weight[92][138],
reservoir_weight[92][139],
reservoir_weight[92][140],
reservoir_weight[92][141],
reservoir_weight[92][142],
reservoir_weight[92][143],
reservoir_weight[92][144],
reservoir_weight[92][145],
reservoir_weight[92][146],
reservoir_weight[92][147],
reservoir_weight[92][148],
reservoir_weight[92][149],
reservoir_weight[92][150],
reservoir_weight[92][151],
reservoir_weight[92][152],
reservoir_weight[92][153],
reservoir_weight[92][154],
reservoir_weight[92][155],
reservoir_weight[92][156],
reservoir_weight[92][157],
reservoir_weight[92][158],
reservoir_weight[92][159],
reservoir_weight[92][160],
reservoir_weight[92][161],
reservoir_weight[92][162],
reservoir_weight[92][163],
reservoir_weight[92][164],
reservoir_weight[92][165],
reservoir_weight[92][166],
reservoir_weight[92][167],
reservoir_weight[92][168],
reservoir_weight[92][169],
reservoir_weight[92][170],
reservoir_weight[92][171],
reservoir_weight[92][172],
reservoir_weight[92][173],
reservoir_weight[92][174],
reservoir_weight[92][175],
reservoir_weight[92][176],
reservoir_weight[92][177],
reservoir_weight[92][178],
reservoir_weight[92][179],
reservoir_weight[92][180],
reservoir_weight[92][181],
reservoir_weight[92][182],
reservoir_weight[92][183],
reservoir_weight[92][184],
reservoir_weight[92][185],
reservoir_weight[92][186],
reservoir_weight[92][187],
reservoir_weight[92][188],
reservoir_weight[92][189],
reservoir_weight[92][190],
reservoir_weight[92][191],
reservoir_weight[92][192],
reservoir_weight[92][193],
reservoir_weight[92][194],
reservoir_weight[92][195],
reservoir_weight[92][196],
reservoir_weight[92][197],
reservoir_weight[92][198],
reservoir_weight[92][199]
},
{reservoir_weight[93][0],
reservoir_weight[93][1],
reservoir_weight[93][2],
reservoir_weight[93][3],
reservoir_weight[93][4],
reservoir_weight[93][5],
reservoir_weight[93][6],
reservoir_weight[93][7],
reservoir_weight[93][8],
reservoir_weight[93][9],
reservoir_weight[93][10],
reservoir_weight[93][11],
reservoir_weight[93][12],
reservoir_weight[93][13],
reservoir_weight[93][14],
reservoir_weight[93][15],
reservoir_weight[93][16],
reservoir_weight[93][17],
reservoir_weight[93][18],
reservoir_weight[93][19],
reservoir_weight[93][20],
reservoir_weight[93][21],
reservoir_weight[93][22],
reservoir_weight[93][23],
reservoir_weight[93][24],
reservoir_weight[93][25],
reservoir_weight[93][26],
reservoir_weight[93][27],
reservoir_weight[93][28],
reservoir_weight[93][29],
reservoir_weight[93][30],
reservoir_weight[93][31],
reservoir_weight[93][32],
reservoir_weight[93][33],
reservoir_weight[93][34],
reservoir_weight[93][35],
reservoir_weight[93][36],
reservoir_weight[93][37],
reservoir_weight[93][38],
reservoir_weight[93][39],
reservoir_weight[93][40],
reservoir_weight[93][41],
reservoir_weight[93][42],
reservoir_weight[93][43],
reservoir_weight[93][44],
reservoir_weight[93][45],
reservoir_weight[93][46],
reservoir_weight[93][47],
reservoir_weight[93][48],
reservoir_weight[93][49],
reservoir_weight[93][50],
reservoir_weight[93][51],
reservoir_weight[93][52],
reservoir_weight[93][53],
reservoir_weight[93][54],
reservoir_weight[93][55],
reservoir_weight[93][56],
reservoir_weight[93][57],
reservoir_weight[93][58],
reservoir_weight[93][59],
reservoir_weight[93][60],
reservoir_weight[93][61],
reservoir_weight[93][62],
reservoir_weight[93][63],
reservoir_weight[93][64],
reservoir_weight[93][65],
reservoir_weight[93][66],
reservoir_weight[93][67],
reservoir_weight[93][68],
reservoir_weight[93][69],
reservoir_weight[93][70],
reservoir_weight[93][71],
reservoir_weight[93][72],
reservoir_weight[93][73],
reservoir_weight[93][74],
reservoir_weight[93][75],
reservoir_weight[93][76],
reservoir_weight[93][77],
reservoir_weight[93][78],
reservoir_weight[93][79],
reservoir_weight[93][80],
reservoir_weight[93][81],
reservoir_weight[93][82],
reservoir_weight[93][83],
reservoir_weight[93][84],
reservoir_weight[93][85],
reservoir_weight[93][86],
reservoir_weight[93][87],
reservoir_weight[93][88],
reservoir_weight[93][89],
reservoir_weight[93][90],
reservoir_weight[93][91],
reservoir_weight[93][92],
reservoir_weight[93][93],
reservoir_weight[93][94],
reservoir_weight[93][95],
reservoir_weight[93][96],
reservoir_weight[93][97],
reservoir_weight[93][98],
reservoir_weight[93][99],
reservoir_weight[93][100],
reservoir_weight[93][101],
reservoir_weight[93][102],
reservoir_weight[93][103],
reservoir_weight[93][104],
reservoir_weight[93][105],
reservoir_weight[93][106],
reservoir_weight[93][107],
reservoir_weight[93][108],
reservoir_weight[93][109],
reservoir_weight[93][110],
reservoir_weight[93][111],
reservoir_weight[93][112],
reservoir_weight[93][113],
reservoir_weight[93][114],
reservoir_weight[93][115],
reservoir_weight[93][116],
reservoir_weight[93][117],
reservoir_weight[93][118],
reservoir_weight[93][119],
reservoir_weight[93][120],
reservoir_weight[93][121],
reservoir_weight[93][122],
reservoir_weight[93][123],
reservoir_weight[93][124],
reservoir_weight[93][125],
reservoir_weight[93][126],
reservoir_weight[93][127],
reservoir_weight[93][128],
reservoir_weight[93][129],
reservoir_weight[93][130],
reservoir_weight[93][131],
reservoir_weight[93][132],
reservoir_weight[93][133],
reservoir_weight[93][134],
reservoir_weight[93][135],
reservoir_weight[93][136],
reservoir_weight[93][137],
reservoir_weight[93][138],
reservoir_weight[93][139],
reservoir_weight[93][140],
reservoir_weight[93][141],
reservoir_weight[93][142],
reservoir_weight[93][143],
reservoir_weight[93][144],
reservoir_weight[93][145],
reservoir_weight[93][146],
reservoir_weight[93][147],
reservoir_weight[93][148],
reservoir_weight[93][149],
reservoir_weight[93][150],
reservoir_weight[93][151],
reservoir_weight[93][152],
reservoir_weight[93][153],
reservoir_weight[93][154],
reservoir_weight[93][155],
reservoir_weight[93][156],
reservoir_weight[93][157],
reservoir_weight[93][158],
reservoir_weight[93][159],
reservoir_weight[93][160],
reservoir_weight[93][161],
reservoir_weight[93][162],
reservoir_weight[93][163],
reservoir_weight[93][164],
reservoir_weight[93][165],
reservoir_weight[93][166],
reservoir_weight[93][167],
reservoir_weight[93][168],
reservoir_weight[93][169],
reservoir_weight[93][170],
reservoir_weight[93][171],
reservoir_weight[93][172],
reservoir_weight[93][173],
reservoir_weight[93][174],
reservoir_weight[93][175],
reservoir_weight[93][176],
reservoir_weight[93][177],
reservoir_weight[93][178],
reservoir_weight[93][179],
reservoir_weight[93][180],
reservoir_weight[93][181],
reservoir_weight[93][182],
reservoir_weight[93][183],
reservoir_weight[93][184],
reservoir_weight[93][185],
reservoir_weight[93][186],
reservoir_weight[93][187],
reservoir_weight[93][188],
reservoir_weight[93][189],
reservoir_weight[93][190],
reservoir_weight[93][191],
reservoir_weight[93][192],
reservoir_weight[93][193],
reservoir_weight[93][194],
reservoir_weight[93][195],
reservoir_weight[93][196],
reservoir_weight[93][197],
reservoir_weight[93][198],
reservoir_weight[93][199]
},
{reservoir_weight[94][0],
reservoir_weight[94][1],
reservoir_weight[94][2],
reservoir_weight[94][3],
reservoir_weight[94][4],
reservoir_weight[94][5],
reservoir_weight[94][6],
reservoir_weight[94][7],
reservoir_weight[94][8],
reservoir_weight[94][9],
reservoir_weight[94][10],
reservoir_weight[94][11],
reservoir_weight[94][12],
reservoir_weight[94][13],
reservoir_weight[94][14],
reservoir_weight[94][15],
reservoir_weight[94][16],
reservoir_weight[94][17],
reservoir_weight[94][18],
reservoir_weight[94][19],
reservoir_weight[94][20],
reservoir_weight[94][21],
reservoir_weight[94][22],
reservoir_weight[94][23],
reservoir_weight[94][24],
reservoir_weight[94][25],
reservoir_weight[94][26],
reservoir_weight[94][27],
reservoir_weight[94][28],
reservoir_weight[94][29],
reservoir_weight[94][30],
reservoir_weight[94][31],
reservoir_weight[94][32],
reservoir_weight[94][33],
reservoir_weight[94][34],
reservoir_weight[94][35],
reservoir_weight[94][36],
reservoir_weight[94][37],
reservoir_weight[94][38],
reservoir_weight[94][39],
reservoir_weight[94][40],
reservoir_weight[94][41],
reservoir_weight[94][42],
reservoir_weight[94][43],
reservoir_weight[94][44],
reservoir_weight[94][45],
reservoir_weight[94][46],
reservoir_weight[94][47],
reservoir_weight[94][48],
reservoir_weight[94][49],
reservoir_weight[94][50],
reservoir_weight[94][51],
reservoir_weight[94][52],
reservoir_weight[94][53],
reservoir_weight[94][54],
reservoir_weight[94][55],
reservoir_weight[94][56],
reservoir_weight[94][57],
reservoir_weight[94][58],
reservoir_weight[94][59],
reservoir_weight[94][60],
reservoir_weight[94][61],
reservoir_weight[94][62],
reservoir_weight[94][63],
reservoir_weight[94][64],
reservoir_weight[94][65],
reservoir_weight[94][66],
reservoir_weight[94][67],
reservoir_weight[94][68],
reservoir_weight[94][69],
reservoir_weight[94][70],
reservoir_weight[94][71],
reservoir_weight[94][72],
reservoir_weight[94][73],
reservoir_weight[94][74],
reservoir_weight[94][75],
reservoir_weight[94][76],
reservoir_weight[94][77],
reservoir_weight[94][78],
reservoir_weight[94][79],
reservoir_weight[94][80],
reservoir_weight[94][81],
reservoir_weight[94][82],
reservoir_weight[94][83],
reservoir_weight[94][84],
reservoir_weight[94][85],
reservoir_weight[94][86],
reservoir_weight[94][87],
reservoir_weight[94][88],
reservoir_weight[94][89],
reservoir_weight[94][90],
reservoir_weight[94][91],
reservoir_weight[94][92],
reservoir_weight[94][93],
reservoir_weight[94][94],
reservoir_weight[94][95],
reservoir_weight[94][96],
reservoir_weight[94][97],
reservoir_weight[94][98],
reservoir_weight[94][99],
reservoir_weight[94][100],
reservoir_weight[94][101],
reservoir_weight[94][102],
reservoir_weight[94][103],
reservoir_weight[94][104],
reservoir_weight[94][105],
reservoir_weight[94][106],
reservoir_weight[94][107],
reservoir_weight[94][108],
reservoir_weight[94][109],
reservoir_weight[94][110],
reservoir_weight[94][111],
reservoir_weight[94][112],
reservoir_weight[94][113],
reservoir_weight[94][114],
reservoir_weight[94][115],
reservoir_weight[94][116],
reservoir_weight[94][117],
reservoir_weight[94][118],
reservoir_weight[94][119],
reservoir_weight[94][120],
reservoir_weight[94][121],
reservoir_weight[94][122],
reservoir_weight[94][123],
reservoir_weight[94][124],
reservoir_weight[94][125],
reservoir_weight[94][126],
reservoir_weight[94][127],
reservoir_weight[94][128],
reservoir_weight[94][129],
reservoir_weight[94][130],
reservoir_weight[94][131],
reservoir_weight[94][132],
reservoir_weight[94][133],
reservoir_weight[94][134],
reservoir_weight[94][135],
reservoir_weight[94][136],
reservoir_weight[94][137],
reservoir_weight[94][138],
reservoir_weight[94][139],
reservoir_weight[94][140],
reservoir_weight[94][141],
reservoir_weight[94][142],
reservoir_weight[94][143],
reservoir_weight[94][144],
reservoir_weight[94][145],
reservoir_weight[94][146],
reservoir_weight[94][147],
reservoir_weight[94][148],
reservoir_weight[94][149],
reservoir_weight[94][150],
reservoir_weight[94][151],
reservoir_weight[94][152],
reservoir_weight[94][153],
reservoir_weight[94][154],
reservoir_weight[94][155],
reservoir_weight[94][156],
reservoir_weight[94][157],
reservoir_weight[94][158],
reservoir_weight[94][159],
reservoir_weight[94][160],
reservoir_weight[94][161],
reservoir_weight[94][162],
reservoir_weight[94][163],
reservoir_weight[94][164],
reservoir_weight[94][165],
reservoir_weight[94][166],
reservoir_weight[94][167],
reservoir_weight[94][168],
reservoir_weight[94][169],
reservoir_weight[94][170],
reservoir_weight[94][171],
reservoir_weight[94][172],
reservoir_weight[94][173],
reservoir_weight[94][174],
reservoir_weight[94][175],
reservoir_weight[94][176],
reservoir_weight[94][177],
reservoir_weight[94][178],
reservoir_weight[94][179],
reservoir_weight[94][180],
reservoir_weight[94][181],
reservoir_weight[94][182],
reservoir_weight[94][183],
reservoir_weight[94][184],
reservoir_weight[94][185],
reservoir_weight[94][186],
reservoir_weight[94][187],
reservoir_weight[94][188],
reservoir_weight[94][189],
reservoir_weight[94][190],
reservoir_weight[94][191],
reservoir_weight[94][192],
reservoir_weight[94][193],
reservoir_weight[94][194],
reservoir_weight[94][195],
reservoir_weight[94][196],
reservoir_weight[94][197],
reservoir_weight[94][198],
reservoir_weight[94][199]
},
{reservoir_weight[95][0],
reservoir_weight[95][1],
reservoir_weight[95][2],
reservoir_weight[95][3],
reservoir_weight[95][4],
reservoir_weight[95][5],
reservoir_weight[95][6],
reservoir_weight[95][7],
reservoir_weight[95][8],
reservoir_weight[95][9],
reservoir_weight[95][10],
reservoir_weight[95][11],
reservoir_weight[95][12],
reservoir_weight[95][13],
reservoir_weight[95][14],
reservoir_weight[95][15],
reservoir_weight[95][16],
reservoir_weight[95][17],
reservoir_weight[95][18],
reservoir_weight[95][19],
reservoir_weight[95][20],
reservoir_weight[95][21],
reservoir_weight[95][22],
reservoir_weight[95][23],
reservoir_weight[95][24],
reservoir_weight[95][25],
reservoir_weight[95][26],
reservoir_weight[95][27],
reservoir_weight[95][28],
reservoir_weight[95][29],
reservoir_weight[95][30],
reservoir_weight[95][31],
reservoir_weight[95][32],
reservoir_weight[95][33],
reservoir_weight[95][34],
reservoir_weight[95][35],
reservoir_weight[95][36],
reservoir_weight[95][37],
reservoir_weight[95][38],
reservoir_weight[95][39],
reservoir_weight[95][40],
reservoir_weight[95][41],
reservoir_weight[95][42],
reservoir_weight[95][43],
reservoir_weight[95][44],
reservoir_weight[95][45],
reservoir_weight[95][46],
reservoir_weight[95][47],
reservoir_weight[95][48],
reservoir_weight[95][49],
reservoir_weight[95][50],
reservoir_weight[95][51],
reservoir_weight[95][52],
reservoir_weight[95][53],
reservoir_weight[95][54],
reservoir_weight[95][55],
reservoir_weight[95][56],
reservoir_weight[95][57],
reservoir_weight[95][58],
reservoir_weight[95][59],
reservoir_weight[95][60],
reservoir_weight[95][61],
reservoir_weight[95][62],
reservoir_weight[95][63],
reservoir_weight[95][64],
reservoir_weight[95][65],
reservoir_weight[95][66],
reservoir_weight[95][67],
reservoir_weight[95][68],
reservoir_weight[95][69],
reservoir_weight[95][70],
reservoir_weight[95][71],
reservoir_weight[95][72],
reservoir_weight[95][73],
reservoir_weight[95][74],
reservoir_weight[95][75],
reservoir_weight[95][76],
reservoir_weight[95][77],
reservoir_weight[95][78],
reservoir_weight[95][79],
reservoir_weight[95][80],
reservoir_weight[95][81],
reservoir_weight[95][82],
reservoir_weight[95][83],
reservoir_weight[95][84],
reservoir_weight[95][85],
reservoir_weight[95][86],
reservoir_weight[95][87],
reservoir_weight[95][88],
reservoir_weight[95][89],
reservoir_weight[95][90],
reservoir_weight[95][91],
reservoir_weight[95][92],
reservoir_weight[95][93],
reservoir_weight[95][94],
reservoir_weight[95][95],
reservoir_weight[95][96],
reservoir_weight[95][97],
reservoir_weight[95][98],
reservoir_weight[95][99],
reservoir_weight[95][100],
reservoir_weight[95][101],
reservoir_weight[95][102],
reservoir_weight[95][103],
reservoir_weight[95][104],
reservoir_weight[95][105],
reservoir_weight[95][106],
reservoir_weight[95][107],
reservoir_weight[95][108],
reservoir_weight[95][109],
reservoir_weight[95][110],
reservoir_weight[95][111],
reservoir_weight[95][112],
reservoir_weight[95][113],
reservoir_weight[95][114],
reservoir_weight[95][115],
reservoir_weight[95][116],
reservoir_weight[95][117],
reservoir_weight[95][118],
reservoir_weight[95][119],
reservoir_weight[95][120],
reservoir_weight[95][121],
reservoir_weight[95][122],
reservoir_weight[95][123],
reservoir_weight[95][124],
reservoir_weight[95][125],
reservoir_weight[95][126],
reservoir_weight[95][127],
reservoir_weight[95][128],
reservoir_weight[95][129],
reservoir_weight[95][130],
reservoir_weight[95][131],
reservoir_weight[95][132],
reservoir_weight[95][133],
reservoir_weight[95][134],
reservoir_weight[95][135],
reservoir_weight[95][136],
reservoir_weight[95][137],
reservoir_weight[95][138],
reservoir_weight[95][139],
reservoir_weight[95][140],
reservoir_weight[95][141],
reservoir_weight[95][142],
reservoir_weight[95][143],
reservoir_weight[95][144],
reservoir_weight[95][145],
reservoir_weight[95][146],
reservoir_weight[95][147],
reservoir_weight[95][148],
reservoir_weight[95][149],
reservoir_weight[95][150],
reservoir_weight[95][151],
reservoir_weight[95][152],
reservoir_weight[95][153],
reservoir_weight[95][154],
reservoir_weight[95][155],
reservoir_weight[95][156],
reservoir_weight[95][157],
reservoir_weight[95][158],
reservoir_weight[95][159],
reservoir_weight[95][160],
reservoir_weight[95][161],
reservoir_weight[95][162],
reservoir_weight[95][163],
reservoir_weight[95][164],
reservoir_weight[95][165],
reservoir_weight[95][166],
reservoir_weight[95][167],
reservoir_weight[95][168],
reservoir_weight[95][169],
reservoir_weight[95][170],
reservoir_weight[95][171],
reservoir_weight[95][172],
reservoir_weight[95][173],
reservoir_weight[95][174],
reservoir_weight[95][175],
reservoir_weight[95][176],
reservoir_weight[95][177],
reservoir_weight[95][178],
reservoir_weight[95][179],
reservoir_weight[95][180],
reservoir_weight[95][181],
reservoir_weight[95][182],
reservoir_weight[95][183],
reservoir_weight[95][184],
reservoir_weight[95][185],
reservoir_weight[95][186],
reservoir_weight[95][187],
reservoir_weight[95][188],
reservoir_weight[95][189],
reservoir_weight[95][190],
reservoir_weight[95][191],
reservoir_weight[95][192],
reservoir_weight[95][193],
reservoir_weight[95][194],
reservoir_weight[95][195],
reservoir_weight[95][196],
reservoir_weight[95][197],
reservoir_weight[95][198],
reservoir_weight[95][199]
},
{reservoir_weight[96][0],
reservoir_weight[96][1],
reservoir_weight[96][2],
reservoir_weight[96][3],
reservoir_weight[96][4],
reservoir_weight[96][5],
reservoir_weight[96][6],
reservoir_weight[96][7],
reservoir_weight[96][8],
reservoir_weight[96][9],
reservoir_weight[96][10],
reservoir_weight[96][11],
reservoir_weight[96][12],
reservoir_weight[96][13],
reservoir_weight[96][14],
reservoir_weight[96][15],
reservoir_weight[96][16],
reservoir_weight[96][17],
reservoir_weight[96][18],
reservoir_weight[96][19],
reservoir_weight[96][20],
reservoir_weight[96][21],
reservoir_weight[96][22],
reservoir_weight[96][23],
reservoir_weight[96][24],
reservoir_weight[96][25],
reservoir_weight[96][26],
reservoir_weight[96][27],
reservoir_weight[96][28],
reservoir_weight[96][29],
reservoir_weight[96][30],
reservoir_weight[96][31],
reservoir_weight[96][32],
reservoir_weight[96][33],
reservoir_weight[96][34],
reservoir_weight[96][35],
reservoir_weight[96][36],
reservoir_weight[96][37],
reservoir_weight[96][38],
reservoir_weight[96][39],
reservoir_weight[96][40],
reservoir_weight[96][41],
reservoir_weight[96][42],
reservoir_weight[96][43],
reservoir_weight[96][44],
reservoir_weight[96][45],
reservoir_weight[96][46],
reservoir_weight[96][47],
reservoir_weight[96][48],
reservoir_weight[96][49],
reservoir_weight[96][50],
reservoir_weight[96][51],
reservoir_weight[96][52],
reservoir_weight[96][53],
reservoir_weight[96][54],
reservoir_weight[96][55],
reservoir_weight[96][56],
reservoir_weight[96][57],
reservoir_weight[96][58],
reservoir_weight[96][59],
reservoir_weight[96][60],
reservoir_weight[96][61],
reservoir_weight[96][62],
reservoir_weight[96][63],
reservoir_weight[96][64],
reservoir_weight[96][65],
reservoir_weight[96][66],
reservoir_weight[96][67],
reservoir_weight[96][68],
reservoir_weight[96][69],
reservoir_weight[96][70],
reservoir_weight[96][71],
reservoir_weight[96][72],
reservoir_weight[96][73],
reservoir_weight[96][74],
reservoir_weight[96][75],
reservoir_weight[96][76],
reservoir_weight[96][77],
reservoir_weight[96][78],
reservoir_weight[96][79],
reservoir_weight[96][80],
reservoir_weight[96][81],
reservoir_weight[96][82],
reservoir_weight[96][83],
reservoir_weight[96][84],
reservoir_weight[96][85],
reservoir_weight[96][86],
reservoir_weight[96][87],
reservoir_weight[96][88],
reservoir_weight[96][89],
reservoir_weight[96][90],
reservoir_weight[96][91],
reservoir_weight[96][92],
reservoir_weight[96][93],
reservoir_weight[96][94],
reservoir_weight[96][95],
reservoir_weight[96][96],
reservoir_weight[96][97],
reservoir_weight[96][98],
reservoir_weight[96][99],
reservoir_weight[96][100],
reservoir_weight[96][101],
reservoir_weight[96][102],
reservoir_weight[96][103],
reservoir_weight[96][104],
reservoir_weight[96][105],
reservoir_weight[96][106],
reservoir_weight[96][107],
reservoir_weight[96][108],
reservoir_weight[96][109],
reservoir_weight[96][110],
reservoir_weight[96][111],
reservoir_weight[96][112],
reservoir_weight[96][113],
reservoir_weight[96][114],
reservoir_weight[96][115],
reservoir_weight[96][116],
reservoir_weight[96][117],
reservoir_weight[96][118],
reservoir_weight[96][119],
reservoir_weight[96][120],
reservoir_weight[96][121],
reservoir_weight[96][122],
reservoir_weight[96][123],
reservoir_weight[96][124],
reservoir_weight[96][125],
reservoir_weight[96][126],
reservoir_weight[96][127],
reservoir_weight[96][128],
reservoir_weight[96][129],
reservoir_weight[96][130],
reservoir_weight[96][131],
reservoir_weight[96][132],
reservoir_weight[96][133],
reservoir_weight[96][134],
reservoir_weight[96][135],
reservoir_weight[96][136],
reservoir_weight[96][137],
reservoir_weight[96][138],
reservoir_weight[96][139],
reservoir_weight[96][140],
reservoir_weight[96][141],
reservoir_weight[96][142],
reservoir_weight[96][143],
reservoir_weight[96][144],
reservoir_weight[96][145],
reservoir_weight[96][146],
reservoir_weight[96][147],
reservoir_weight[96][148],
reservoir_weight[96][149],
reservoir_weight[96][150],
reservoir_weight[96][151],
reservoir_weight[96][152],
reservoir_weight[96][153],
reservoir_weight[96][154],
reservoir_weight[96][155],
reservoir_weight[96][156],
reservoir_weight[96][157],
reservoir_weight[96][158],
reservoir_weight[96][159],
reservoir_weight[96][160],
reservoir_weight[96][161],
reservoir_weight[96][162],
reservoir_weight[96][163],
reservoir_weight[96][164],
reservoir_weight[96][165],
reservoir_weight[96][166],
reservoir_weight[96][167],
reservoir_weight[96][168],
reservoir_weight[96][169],
reservoir_weight[96][170],
reservoir_weight[96][171],
reservoir_weight[96][172],
reservoir_weight[96][173],
reservoir_weight[96][174],
reservoir_weight[96][175],
reservoir_weight[96][176],
reservoir_weight[96][177],
reservoir_weight[96][178],
reservoir_weight[96][179],
reservoir_weight[96][180],
reservoir_weight[96][181],
reservoir_weight[96][182],
reservoir_weight[96][183],
reservoir_weight[96][184],
reservoir_weight[96][185],
reservoir_weight[96][186],
reservoir_weight[96][187],
reservoir_weight[96][188],
reservoir_weight[96][189],
reservoir_weight[96][190],
reservoir_weight[96][191],
reservoir_weight[96][192],
reservoir_weight[96][193],
reservoir_weight[96][194],
reservoir_weight[96][195],
reservoir_weight[96][196],
reservoir_weight[96][197],
reservoir_weight[96][198],
reservoir_weight[96][199]
},
{reservoir_weight[97][0],
reservoir_weight[97][1],
reservoir_weight[97][2],
reservoir_weight[97][3],
reservoir_weight[97][4],
reservoir_weight[97][5],
reservoir_weight[97][6],
reservoir_weight[97][7],
reservoir_weight[97][8],
reservoir_weight[97][9],
reservoir_weight[97][10],
reservoir_weight[97][11],
reservoir_weight[97][12],
reservoir_weight[97][13],
reservoir_weight[97][14],
reservoir_weight[97][15],
reservoir_weight[97][16],
reservoir_weight[97][17],
reservoir_weight[97][18],
reservoir_weight[97][19],
reservoir_weight[97][20],
reservoir_weight[97][21],
reservoir_weight[97][22],
reservoir_weight[97][23],
reservoir_weight[97][24],
reservoir_weight[97][25],
reservoir_weight[97][26],
reservoir_weight[97][27],
reservoir_weight[97][28],
reservoir_weight[97][29],
reservoir_weight[97][30],
reservoir_weight[97][31],
reservoir_weight[97][32],
reservoir_weight[97][33],
reservoir_weight[97][34],
reservoir_weight[97][35],
reservoir_weight[97][36],
reservoir_weight[97][37],
reservoir_weight[97][38],
reservoir_weight[97][39],
reservoir_weight[97][40],
reservoir_weight[97][41],
reservoir_weight[97][42],
reservoir_weight[97][43],
reservoir_weight[97][44],
reservoir_weight[97][45],
reservoir_weight[97][46],
reservoir_weight[97][47],
reservoir_weight[97][48],
reservoir_weight[97][49],
reservoir_weight[97][50],
reservoir_weight[97][51],
reservoir_weight[97][52],
reservoir_weight[97][53],
reservoir_weight[97][54],
reservoir_weight[97][55],
reservoir_weight[97][56],
reservoir_weight[97][57],
reservoir_weight[97][58],
reservoir_weight[97][59],
reservoir_weight[97][60],
reservoir_weight[97][61],
reservoir_weight[97][62],
reservoir_weight[97][63],
reservoir_weight[97][64],
reservoir_weight[97][65],
reservoir_weight[97][66],
reservoir_weight[97][67],
reservoir_weight[97][68],
reservoir_weight[97][69],
reservoir_weight[97][70],
reservoir_weight[97][71],
reservoir_weight[97][72],
reservoir_weight[97][73],
reservoir_weight[97][74],
reservoir_weight[97][75],
reservoir_weight[97][76],
reservoir_weight[97][77],
reservoir_weight[97][78],
reservoir_weight[97][79],
reservoir_weight[97][80],
reservoir_weight[97][81],
reservoir_weight[97][82],
reservoir_weight[97][83],
reservoir_weight[97][84],
reservoir_weight[97][85],
reservoir_weight[97][86],
reservoir_weight[97][87],
reservoir_weight[97][88],
reservoir_weight[97][89],
reservoir_weight[97][90],
reservoir_weight[97][91],
reservoir_weight[97][92],
reservoir_weight[97][93],
reservoir_weight[97][94],
reservoir_weight[97][95],
reservoir_weight[97][96],
reservoir_weight[97][97],
reservoir_weight[97][98],
reservoir_weight[97][99],
reservoir_weight[97][100],
reservoir_weight[97][101],
reservoir_weight[97][102],
reservoir_weight[97][103],
reservoir_weight[97][104],
reservoir_weight[97][105],
reservoir_weight[97][106],
reservoir_weight[97][107],
reservoir_weight[97][108],
reservoir_weight[97][109],
reservoir_weight[97][110],
reservoir_weight[97][111],
reservoir_weight[97][112],
reservoir_weight[97][113],
reservoir_weight[97][114],
reservoir_weight[97][115],
reservoir_weight[97][116],
reservoir_weight[97][117],
reservoir_weight[97][118],
reservoir_weight[97][119],
reservoir_weight[97][120],
reservoir_weight[97][121],
reservoir_weight[97][122],
reservoir_weight[97][123],
reservoir_weight[97][124],
reservoir_weight[97][125],
reservoir_weight[97][126],
reservoir_weight[97][127],
reservoir_weight[97][128],
reservoir_weight[97][129],
reservoir_weight[97][130],
reservoir_weight[97][131],
reservoir_weight[97][132],
reservoir_weight[97][133],
reservoir_weight[97][134],
reservoir_weight[97][135],
reservoir_weight[97][136],
reservoir_weight[97][137],
reservoir_weight[97][138],
reservoir_weight[97][139],
reservoir_weight[97][140],
reservoir_weight[97][141],
reservoir_weight[97][142],
reservoir_weight[97][143],
reservoir_weight[97][144],
reservoir_weight[97][145],
reservoir_weight[97][146],
reservoir_weight[97][147],
reservoir_weight[97][148],
reservoir_weight[97][149],
reservoir_weight[97][150],
reservoir_weight[97][151],
reservoir_weight[97][152],
reservoir_weight[97][153],
reservoir_weight[97][154],
reservoir_weight[97][155],
reservoir_weight[97][156],
reservoir_weight[97][157],
reservoir_weight[97][158],
reservoir_weight[97][159],
reservoir_weight[97][160],
reservoir_weight[97][161],
reservoir_weight[97][162],
reservoir_weight[97][163],
reservoir_weight[97][164],
reservoir_weight[97][165],
reservoir_weight[97][166],
reservoir_weight[97][167],
reservoir_weight[97][168],
reservoir_weight[97][169],
reservoir_weight[97][170],
reservoir_weight[97][171],
reservoir_weight[97][172],
reservoir_weight[97][173],
reservoir_weight[97][174],
reservoir_weight[97][175],
reservoir_weight[97][176],
reservoir_weight[97][177],
reservoir_weight[97][178],
reservoir_weight[97][179],
reservoir_weight[97][180],
reservoir_weight[97][181],
reservoir_weight[97][182],
reservoir_weight[97][183],
reservoir_weight[97][184],
reservoir_weight[97][185],
reservoir_weight[97][186],
reservoir_weight[97][187],
reservoir_weight[97][188],
reservoir_weight[97][189],
reservoir_weight[97][190],
reservoir_weight[97][191],
reservoir_weight[97][192],
reservoir_weight[97][193],
reservoir_weight[97][194],
reservoir_weight[97][195],
reservoir_weight[97][196],
reservoir_weight[97][197],
reservoir_weight[97][198],
reservoir_weight[97][199]
},
{reservoir_weight[98][0],
reservoir_weight[98][1],
reservoir_weight[98][2],
reservoir_weight[98][3],
reservoir_weight[98][4],
reservoir_weight[98][5],
reservoir_weight[98][6],
reservoir_weight[98][7],
reservoir_weight[98][8],
reservoir_weight[98][9],
reservoir_weight[98][10],
reservoir_weight[98][11],
reservoir_weight[98][12],
reservoir_weight[98][13],
reservoir_weight[98][14],
reservoir_weight[98][15],
reservoir_weight[98][16],
reservoir_weight[98][17],
reservoir_weight[98][18],
reservoir_weight[98][19],
reservoir_weight[98][20],
reservoir_weight[98][21],
reservoir_weight[98][22],
reservoir_weight[98][23],
reservoir_weight[98][24],
reservoir_weight[98][25],
reservoir_weight[98][26],
reservoir_weight[98][27],
reservoir_weight[98][28],
reservoir_weight[98][29],
reservoir_weight[98][30],
reservoir_weight[98][31],
reservoir_weight[98][32],
reservoir_weight[98][33],
reservoir_weight[98][34],
reservoir_weight[98][35],
reservoir_weight[98][36],
reservoir_weight[98][37],
reservoir_weight[98][38],
reservoir_weight[98][39],
reservoir_weight[98][40],
reservoir_weight[98][41],
reservoir_weight[98][42],
reservoir_weight[98][43],
reservoir_weight[98][44],
reservoir_weight[98][45],
reservoir_weight[98][46],
reservoir_weight[98][47],
reservoir_weight[98][48],
reservoir_weight[98][49],
reservoir_weight[98][50],
reservoir_weight[98][51],
reservoir_weight[98][52],
reservoir_weight[98][53],
reservoir_weight[98][54],
reservoir_weight[98][55],
reservoir_weight[98][56],
reservoir_weight[98][57],
reservoir_weight[98][58],
reservoir_weight[98][59],
reservoir_weight[98][60],
reservoir_weight[98][61],
reservoir_weight[98][62],
reservoir_weight[98][63],
reservoir_weight[98][64],
reservoir_weight[98][65],
reservoir_weight[98][66],
reservoir_weight[98][67],
reservoir_weight[98][68],
reservoir_weight[98][69],
reservoir_weight[98][70],
reservoir_weight[98][71],
reservoir_weight[98][72],
reservoir_weight[98][73],
reservoir_weight[98][74],
reservoir_weight[98][75],
reservoir_weight[98][76],
reservoir_weight[98][77],
reservoir_weight[98][78],
reservoir_weight[98][79],
reservoir_weight[98][80],
reservoir_weight[98][81],
reservoir_weight[98][82],
reservoir_weight[98][83],
reservoir_weight[98][84],
reservoir_weight[98][85],
reservoir_weight[98][86],
reservoir_weight[98][87],
reservoir_weight[98][88],
reservoir_weight[98][89],
reservoir_weight[98][90],
reservoir_weight[98][91],
reservoir_weight[98][92],
reservoir_weight[98][93],
reservoir_weight[98][94],
reservoir_weight[98][95],
reservoir_weight[98][96],
reservoir_weight[98][97],
reservoir_weight[98][98],
reservoir_weight[98][99],
reservoir_weight[98][100],
reservoir_weight[98][101],
reservoir_weight[98][102],
reservoir_weight[98][103],
reservoir_weight[98][104],
reservoir_weight[98][105],
reservoir_weight[98][106],
reservoir_weight[98][107],
reservoir_weight[98][108],
reservoir_weight[98][109],
reservoir_weight[98][110],
reservoir_weight[98][111],
reservoir_weight[98][112],
reservoir_weight[98][113],
reservoir_weight[98][114],
reservoir_weight[98][115],
reservoir_weight[98][116],
reservoir_weight[98][117],
reservoir_weight[98][118],
reservoir_weight[98][119],
reservoir_weight[98][120],
reservoir_weight[98][121],
reservoir_weight[98][122],
reservoir_weight[98][123],
reservoir_weight[98][124],
reservoir_weight[98][125],
reservoir_weight[98][126],
reservoir_weight[98][127],
reservoir_weight[98][128],
reservoir_weight[98][129],
reservoir_weight[98][130],
reservoir_weight[98][131],
reservoir_weight[98][132],
reservoir_weight[98][133],
reservoir_weight[98][134],
reservoir_weight[98][135],
reservoir_weight[98][136],
reservoir_weight[98][137],
reservoir_weight[98][138],
reservoir_weight[98][139],
reservoir_weight[98][140],
reservoir_weight[98][141],
reservoir_weight[98][142],
reservoir_weight[98][143],
reservoir_weight[98][144],
reservoir_weight[98][145],
reservoir_weight[98][146],
reservoir_weight[98][147],
reservoir_weight[98][148],
reservoir_weight[98][149],
reservoir_weight[98][150],
reservoir_weight[98][151],
reservoir_weight[98][152],
reservoir_weight[98][153],
reservoir_weight[98][154],
reservoir_weight[98][155],
reservoir_weight[98][156],
reservoir_weight[98][157],
reservoir_weight[98][158],
reservoir_weight[98][159],
reservoir_weight[98][160],
reservoir_weight[98][161],
reservoir_weight[98][162],
reservoir_weight[98][163],
reservoir_weight[98][164],
reservoir_weight[98][165],
reservoir_weight[98][166],
reservoir_weight[98][167],
reservoir_weight[98][168],
reservoir_weight[98][169],
reservoir_weight[98][170],
reservoir_weight[98][171],
reservoir_weight[98][172],
reservoir_weight[98][173],
reservoir_weight[98][174],
reservoir_weight[98][175],
reservoir_weight[98][176],
reservoir_weight[98][177],
reservoir_weight[98][178],
reservoir_weight[98][179],
reservoir_weight[98][180],
reservoir_weight[98][181],
reservoir_weight[98][182],
reservoir_weight[98][183],
reservoir_weight[98][184],
reservoir_weight[98][185],
reservoir_weight[98][186],
reservoir_weight[98][187],
reservoir_weight[98][188],
reservoir_weight[98][189],
reservoir_weight[98][190],
reservoir_weight[98][191],
reservoir_weight[98][192],
reservoir_weight[98][193],
reservoir_weight[98][194],
reservoir_weight[98][195],
reservoir_weight[98][196],
reservoir_weight[98][197],
reservoir_weight[98][198],
reservoir_weight[98][199]
},
{reservoir_weight[99][0],
reservoir_weight[99][1],
reservoir_weight[99][2],
reservoir_weight[99][3],
reservoir_weight[99][4],
reservoir_weight[99][5],
reservoir_weight[99][6],
reservoir_weight[99][7],
reservoir_weight[99][8],
reservoir_weight[99][9],
reservoir_weight[99][10],
reservoir_weight[99][11],
reservoir_weight[99][12],
reservoir_weight[99][13],
reservoir_weight[99][14],
reservoir_weight[99][15],
reservoir_weight[99][16],
reservoir_weight[99][17],
reservoir_weight[99][18],
reservoir_weight[99][19],
reservoir_weight[99][20],
reservoir_weight[99][21],
reservoir_weight[99][22],
reservoir_weight[99][23],
reservoir_weight[99][24],
reservoir_weight[99][25],
reservoir_weight[99][26],
reservoir_weight[99][27],
reservoir_weight[99][28],
reservoir_weight[99][29],
reservoir_weight[99][30],
reservoir_weight[99][31],
reservoir_weight[99][32],
reservoir_weight[99][33],
reservoir_weight[99][34],
reservoir_weight[99][35],
reservoir_weight[99][36],
reservoir_weight[99][37],
reservoir_weight[99][38],
reservoir_weight[99][39],
reservoir_weight[99][40],
reservoir_weight[99][41],
reservoir_weight[99][42],
reservoir_weight[99][43],
reservoir_weight[99][44],
reservoir_weight[99][45],
reservoir_weight[99][46],
reservoir_weight[99][47],
reservoir_weight[99][48],
reservoir_weight[99][49],
reservoir_weight[99][50],
reservoir_weight[99][51],
reservoir_weight[99][52],
reservoir_weight[99][53],
reservoir_weight[99][54],
reservoir_weight[99][55],
reservoir_weight[99][56],
reservoir_weight[99][57],
reservoir_weight[99][58],
reservoir_weight[99][59],
reservoir_weight[99][60],
reservoir_weight[99][61],
reservoir_weight[99][62],
reservoir_weight[99][63],
reservoir_weight[99][64],
reservoir_weight[99][65],
reservoir_weight[99][66],
reservoir_weight[99][67],
reservoir_weight[99][68],
reservoir_weight[99][69],
reservoir_weight[99][70],
reservoir_weight[99][71],
reservoir_weight[99][72],
reservoir_weight[99][73],
reservoir_weight[99][74],
reservoir_weight[99][75],
reservoir_weight[99][76],
reservoir_weight[99][77],
reservoir_weight[99][78],
reservoir_weight[99][79],
reservoir_weight[99][80],
reservoir_weight[99][81],
reservoir_weight[99][82],
reservoir_weight[99][83],
reservoir_weight[99][84],
reservoir_weight[99][85],
reservoir_weight[99][86],
reservoir_weight[99][87],
reservoir_weight[99][88],
reservoir_weight[99][89],
reservoir_weight[99][90],
reservoir_weight[99][91],
reservoir_weight[99][92],
reservoir_weight[99][93],
reservoir_weight[99][94],
reservoir_weight[99][95],
reservoir_weight[99][96],
reservoir_weight[99][97],
reservoir_weight[99][98],
reservoir_weight[99][99],
reservoir_weight[99][100],
reservoir_weight[99][101],
reservoir_weight[99][102],
reservoir_weight[99][103],
reservoir_weight[99][104],
reservoir_weight[99][105],
reservoir_weight[99][106],
reservoir_weight[99][107],
reservoir_weight[99][108],
reservoir_weight[99][109],
reservoir_weight[99][110],
reservoir_weight[99][111],
reservoir_weight[99][112],
reservoir_weight[99][113],
reservoir_weight[99][114],
reservoir_weight[99][115],
reservoir_weight[99][116],
reservoir_weight[99][117],
reservoir_weight[99][118],
reservoir_weight[99][119],
reservoir_weight[99][120],
reservoir_weight[99][121],
reservoir_weight[99][122],
reservoir_weight[99][123],
reservoir_weight[99][124],
reservoir_weight[99][125],
reservoir_weight[99][126],
reservoir_weight[99][127],
reservoir_weight[99][128],
reservoir_weight[99][129],
reservoir_weight[99][130],
reservoir_weight[99][131],
reservoir_weight[99][132],
reservoir_weight[99][133],
reservoir_weight[99][134],
reservoir_weight[99][135],
reservoir_weight[99][136],
reservoir_weight[99][137],
reservoir_weight[99][138],
reservoir_weight[99][139],
reservoir_weight[99][140],
reservoir_weight[99][141],
reservoir_weight[99][142],
reservoir_weight[99][143],
reservoir_weight[99][144],
reservoir_weight[99][145],
reservoir_weight[99][146],
reservoir_weight[99][147],
reservoir_weight[99][148],
reservoir_weight[99][149],
reservoir_weight[99][150],
reservoir_weight[99][151],
reservoir_weight[99][152],
reservoir_weight[99][153],
reservoir_weight[99][154],
reservoir_weight[99][155],
reservoir_weight[99][156],
reservoir_weight[99][157],
reservoir_weight[99][158],
reservoir_weight[99][159],
reservoir_weight[99][160],
reservoir_weight[99][161],
reservoir_weight[99][162],
reservoir_weight[99][163],
reservoir_weight[99][164],
reservoir_weight[99][165],
reservoir_weight[99][166],
reservoir_weight[99][167],
reservoir_weight[99][168],
reservoir_weight[99][169],
reservoir_weight[99][170],
reservoir_weight[99][171],
reservoir_weight[99][172],
reservoir_weight[99][173],
reservoir_weight[99][174],
reservoir_weight[99][175],
reservoir_weight[99][176],
reservoir_weight[99][177],
reservoir_weight[99][178],
reservoir_weight[99][179],
reservoir_weight[99][180],
reservoir_weight[99][181],
reservoir_weight[99][182],
reservoir_weight[99][183],
reservoir_weight[99][184],
reservoir_weight[99][185],
reservoir_weight[99][186],
reservoir_weight[99][187],
reservoir_weight[99][188],
reservoir_weight[99][189],
reservoir_weight[99][190],
reservoir_weight[99][191],
reservoir_weight[99][192],
reservoir_weight[99][193],
reservoir_weight[99][194],
reservoir_weight[99][195],
reservoir_weight[99][196],
reservoir_weight[99][197],
reservoir_weight[99][198],
reservoir_weight[99][199]
},
{reservoir_weight[100][0],
reservoir_weight[100][1],
reservoir_weight[100][2],
reservoir_weight[100][3],
reservoir_weight[100][4],
reservoir_weight[100][5],
reservoir_weight[100][6],
reservoir_weight[100][7],
reservoir_weight[100][8],
reservoir_weight[100][9],
reservoir_weight[100][10],
reservoir_weight[100][11],
reservoir_weight[100][12],
reservoir_weight[100][13],
reservoir_weight[100][14],
reservoir_weight[100][15],
reservoir_weight[100][16],
reservoir_weight[100][17],
reservoir_weight[100][18],
reservoir_weight[100][19],
reservoir_weight[100][20],
reservoir_weight[100][21],
reservoir_weight[100][22],
reservoir_weight[100][23],
reservoir_weight[100][24],
reservoir_weight[100][25],
reservoir_weight[100][26],
reservoir_weight[100][27],
reservoir_weight[100][28],
reservoir_weight[100][29],
reservoir_weight[100][30],
reservoir_weight[100][31],
reservoir_weight[100][32],
reservoir_weight[100][33],
reservoir_weight[100][34],
reservoir_weight[100][35],
reservoir_weight[100][36],
reservoir_weight[100][37],
reservoir_weight[100][38],
reservoir_weight[100][39],
reservoir_weight[100][40],
reservoir_weight[100][41],
reservoir_weight[100][42],
reservoir_weight[100][43],
reservoir_weight[100][44],
reservoir_weight[100][45],
reservoir_weight[100][46],
reservoir_weight[100][47],
reservoir_weight[100][48],
reservoir_weight[100][49],
reservoir_weight[100][50],
reservoir_weight[100][51],
reservoir_weight[100][52],
reservoir_weight[100][53],
reservoir_weight[100][54],
reservoir_weight[100][55],
reservoir_weight[100][56],
reservoir_weight[100][57],
reservoir_weight[100][58],
reservoir_weight[100][59],
reservoir_weight[100][60],
reservoir_weight[100][61],
reservoir_weight[100][62],
reservoir_weight[100][63],
reservoir_weight[100][64],
reservoir_weight[100][65],
reservoir_weight[100][66],
reservoir_weight[100][67],
reservoir_weight[100][68],
reservoir_weight[100][69],
reservoir_weight[100][70],
reservoir_weight[100][71],
reservoir_weight[100][72],
reservoir_weight[100][73],
reservoir_weight[100][74],
reservoir_weight[100][75],
reservoir_weight[100][76],
reservoir_weight[100][77],
reservoir_weight[100][78],
reservoir_weight[100][79],
reservoir_weight[100][80],
reservoir_weight[100][81],
reservoir_weight[100][82],
reservoir_weight[100][83],
reservoir_weight[100][84],
reservoir_weight[100][85],
reservoir_weight[100][86],
reservoir_weight[100][87],
reservoir_weight[100][88],
reservoir_weight[100][89],
reservoir_weight[100][90],
reservoir_weight[100][91],
reservoir_weight[100][92],
reservoir_weight[100][93],
reservoir_weight[100][94],
reservoir_weight[100][95],
reservoir_weight[100][96],
reservoir_weight[100][97],
reservoir_weight[100][98],
reservoir_weight[100][99],
reservoir_weight[100][100],
reservoir_weight[100][101],
reservoir_weight[100][102],
reservoir_weight[100][103],
reservoir_weight[100][104],
reservoir_weight[100][105],
reservoir_weight[100][106],
reservoir_weight[100][107],
reservoir_weight[100][108],
reservoir_weight[100][109],
reservoir_weight[100][110],
reservoir_weight[100][111],
reservoir_weight[100][112],
reservoir_weight[100][113],
reservoir_weight[100][114],
reservoir_weight[100][115],
reservoir_weight[100][116],
reservoir_weight[100][117],
reservoir_weight[100][118],
reservoir_weight[100][119],
reservoir_weight[100][120],
reservoir_weight[100][121],
reservoir_weight[100][122],
reservoir_weight[100][123],
reservoir_weight[100][124],
reservoir_weight[100][125],
reservoir_weight[100][126],
reservoir_weight[100][127],
reservoir_weight[100][128],
reservoir_weight[100][129],
reservoir_weight[100][130],
reservoir_weight[100][131],
reservoir_weight[100][132],
reservoir_weight[100][133],
reservoir_weight[100][134],
reservoir_weight[100][135],
reservoir_weight[100][136],
reservoir_weight[100][137],
reservoir_weight[100][138],
reservoir_weight[100][139],
reservoir_weight[100][140],
reservoir_weight[100][141],
reservoir_weight[100][142],
reservoir_weight[100][143],
reservoir_weight[100][144],
reservoir_weight[100][145],
reservoir_weight[100][146],
reservoir_weight[100][147],
reservoir_weight[100][148],
reservoir_weight[100][149],
reservoir_weight[100][150],
reservoir_weight[100][151],
reservoir_weight[100][152],
reservoir_weight[100][153],
reservoir_weight[100][154],
reservoir_weight[100][155],
reservoir_weight[100][156],
reservoir_weight[100][157],
reservoir_weight[100][158],
reservoir_weight[100][159],
reservoir_weight[100][160],
reservoir_weight[100][161],
reservoir_weight[100][162],
reservoir_weight[100][163],
reservoir_weight[100][164],
reservoir_weight[100][165],
reservoir_weight[100][166],
reservoir_weight[100][167],
reservoir_weight[100][168],
reservoir_weight[100][169],
reservoir_weight[100][170],
reservoir_weight[100][171],
reservoir_weight[100][172],
reservoir_weight[100][173],
reservoir_weight[100][174],
reservoir_weight[100][175],
reservoir_weight[100][176],
reservoir_weight[100][177],
reservoir_weight[100][178],
reservoir_weight[100][179],
reservoir_weight[100][180],
reservoir_weight[100][181],
reservoir_weight[100][182],
reservoir_weight[100][183],
reservoir_weight[100][184],
reservoir_weight[100][185],
reservoir_weight[100][186],
reservoir_weight[100][187],
reservoir_weight[100][188],
reservoir_weight[100][189],
reservoir_weight[100][190],
reservoir_weight[100][191],
reservoir_weight[100][192],
reservoir_weight[100][193],
reservoir_weight[100][194],
reservoir_weight[100][195],
reservoir_weight[100][196],
reservoir_weight[100][197],
reservoir_weight[100][198],
reservoir_weight[100][199]
},
{reservoir_weight[101][0],
reservoir_weight[101][1],
reservoir_weight[101][2],
reservoir_weight[101][3],
reservoir_weight[101][4],
reservoir_weight[101][5],
reservoir_weight[101][6],
reservoir_weight[101][7],
reservoir_weight[101][8],
reservoir_weight[101][9],
reservoir_weight[101][10],
reservoir_weight[101][11],
reservoir_weight[101][12],
reservoir_weight[101][13],
reservoir_weight[101][14],
reservoir_weight[101][15],
reservoir_weight[101][16],
reservoir_weight[101][17],
reservoir_weight[101][18],
reservoir_weight[101][19],
reservoir_weight[101][20],
reservoir_weight[101][21],
reservoir_weight[101][22],
reservoir_weight[101][23],
reservoir_weight[101][24],
reservoir_weight[101][25],
reservoir_weight[101][26],
reservoir_weight[101][27],
reservoir_weight[101][28],
reservoir_weight[101][29],
reservoir_weight[101][30],
reservoir_weight[101][31],
reservoir_weight[101][32],
reservoir_weight[101][33],
reservoir_weight[101][34],
reservoir_weight[101][35],
reservoir_weight[101][36],
reservoir_weight[101][37],
reservoir_weight[101][38],
reservoir_weight[101][39],
reservoir_weight[101][40],
reservoir_weight[101][41],
reservoir_weight[101][42],
reservoir_weight[101][43],
reservoir_weight[101][44],
reservoir_weight[101][45],
reservoir_weight[101][46],
reservoir_weight[101][47],
reservoir_weight[101][48],
reservoir_weight[101][49],
reservoir_weight[101][50],
reservoir_weight[101][51],
reservoir_weight[101][52],
reservoir_weight[101][53],
reservoir_weight[101][54],
reservoir_weight[101][55],
reservoir_weight[101][56],
reservoir_weight[101][57],
reservoir_weight[101][58],
reservoir_weight[101][59],
reservoir_weight[101][60],
reservoir_weight[101][61],
reservoir_weight[101][62],
reservoir_weight[101][63],
reservoir_weight[101][64],
reservoir_weight[101][65],
reservoir_weight[101][66],
reservoir_weight[101][67],
reservoir_weight[101][68],
reservoir_weight[101][69],
reservoir_weight[101][70],
reservoir_weight[101][71],
reservoir_weight[101][72],
reservoir_weight[101][73],
reservoir_weight[101][74],
reservoir_weight[101][75],
reservoir_weight[101][76],
reservoir_weight[101][77],
reservoir_weight[101][78],
reservoir_weight[101][79],
reservoir_weight[101][80],
reservoir_weight[101][81],
reservoir_weight[101][82],
reservoir_weight[101][83],
reservoir_weight[101][84],
reservoir_weight[101][85],
reservoir_weight[101][86],
reservoir_weight[101][87],
reservoir_weight[101][88],
reservoir_weight[101][89],
reservoir_weight[101][90],
reservoir_weight[101][91],
reservoir_weight[101][92],
reservoir_weight[101][93],
reservoir_weight[101][94],
reservoir_weight[101][95],
reservoir_weight[101][96],
reservoir_weight[101][97],
reservoir_weight[101][98],
reservoir_weight[101][99],
reservoir_weight[101][100],
reservoir_weight[101][101],
reservoir_weight[101][102],
reservoir_weight[101][103],
reservoir_weight[101][104],
reservoir_weight[101][105],
reservoir_weight[101][106],
reservoir_weight[101][107],
reservoir_weight[101][108],
reservoir_weight[101][109],
reservoir_weight[101][110],
reservoir_weight[101][111],
reservoir_weight[101][112],
reservoir_weight[101][113],
reservoir_weight[101][114],
reservoir_weight[101][115],
reservoir_weight[101][116],
reservoir_weight[101][117],
reservoir_weight[101][118],
reservoir_weight[101][119],
reservoir_weight[101][120],
reservoir_weight[101][121],
reservoir_weight[101][122],
reservoir_weight[101][123],
reservoir_weight[101][124],
reservoir_weight[101][125],
reservoir_weight[101][126],
reservoir_weight[101][127],
reservoir_weight[101][128],
reservoir_weight[101][129],
reservoir_weight[101][130],
reservoir_weight[101][131],
reservoir_weight[101][132],
reservoir_weight[101][133],
reservoir_weight[101][134],
reservoir_weight[101][135],
reservoir_weight[101][136],
reservoir_weight[101][137],
reservoir_weight[101][138],
reservoir_weight[101][139],
reservoir_weight[101][140],
reservoir_weight[101][141],
reservoir_weight[101][142],
reservoir_weight[101][143],
reservoir_weight[101][144],
reservoir_weight[101][145],
reservoir_weight[101][146],
reservoir_weight[101][147],
reservoir_weight[101][148],
reservoir_weight[101][149],
reservoir_weight[101][150],
reservoir_weight[101][151],
reservoir_weight[101][152],
reservoir_weight[101][153],
reservoir_weight[101][154],
reservoir_weight[101][155],
reservoir_weight[101][156],
reservoir_weight[101][157],
reservoir_weight[101][158],
reservoir_weight[101][159],
reservoir_weight[101][160],
reservoir_weight[101][161],
reservoir_weight[101][162],
reservoir_weight[101][163],
reservoir_weight[101][164],
reservoir_weight[101][165],
reservoir_weight[101][166],
reservoir_weight[101][167],
reservoir_weight[101][168],
reservoir_weight[101][169],
reservoir_weight[101][170],
reservoir_weight[101][171],
reservoir_weight[101][172],
reservoir_weight[101][173],
reservoir_weight[101][174],
reservoir_weight[101][175],
reservoir_weight[101][176],
reservoir_weight[101][177],
reservoir_weight[101][178],
reservoir_weight[101][179],
reservoir_weight[101][180],
reservoir_weight[101][181],
reservoir_weight[101][182],
reservoir_weight[101][183],
reservoir_weight[101][184],
reservoir_weight[101][185],
reservoir_weight[101][186],
reservoir_weight[101][187],
reservoir_weight[101][188],
reservoir_weight[101][189],
reservoir_weight[101][190],
reservoir_weight[101][191],
reservoir_weight[101][192],
reservoir_weight[101][193],
reservoir_weight[101][194],
reservoir_weight[101][195],
reservoir_weight[101][196],
reservoir_weight[101][197],
reservoir_weight[101][198],
reservoir_weight[101][199]
},
{reservoir_weight[102][0],
reservoir_weight[102][1],
reservoir_weight[102][2],
reservoir_weight[102][3],
reservoir_weight[102][4],
reservoir_weight[102][5],
reservoir_weight[102][6],
reservoir_weight[102][7],
reservoir_weight[102][8],
reservoir_weight[102][9],
reservoir_weight[102][10],
reservoir_weight[102][11],
reservoir_weight[102][12],
reservoir_weight[102][13],
reservoir_weight[102][14],
reservoir_weight[102][15],
reservoir_weight[102][16],
reservoir_weight[102][17],
reservoir_weight[102][18],
reservoir_weight[102][19],
reservoir_weight[102][20],
reservoir_weight[102][21],
reservoir_weight[102][22],
reservoir_weight[102][23],
reservoir_weight[102][24],
reservoir_weight[102][25],
reservoir_weight[102][26],
reservoir_weight[102][27],
reservoir_weight[102][28],
reservoir_weight[102][29],
reservoir_weight[102][30],
reservoir_weight[102][31],
reservoir_weight[102][32],
reservoir_weight[102][33],
reservoir_weight[102][34],
reservoir_weight[102][35],
reservoir_weight[102][36],
reservoir_weight[102][37],
reservoir_weight[102][38],
reservoir_weight[102][39],
reservoir_weight[102][40],
reservoir_weight[102][41],
reservoir_weight[102][42],
reservoir_weight[102][43],
reservoir_weight[102][44],
reservoir_weight[102][45],
reservoir_weight[102][46],
reservoir_weight[102][47],
reservoir_weight[102][48],
reservoir_weight[102][49],
reservoir_weight[102][50],
reservoir_weight[102][51],
reservoir_weight[102][52],
reservoir_weight[102][53],
reservoir_weight[102][54],
reservoir_weight[102][55],
reservoir_weight[102][56],
reservoir_weight[102][57],
reservoir_weight[102][58],
reservoir_weight[102][59],
reservoir_weight[102][60],
reservoir_weight[102][61],
reservoir_weight[102][62],
reservoir_weight[102][63],
reservoir_weight[102][64],
reservoir_weight[102][65],
reservoir_weight[102][66],
reservoir_weight[102][67],
reservoir_weight[102][68],
reservoir_weight[102][69],
reservoir_weight[102][70],
reservoir_weight[102][71],
reservoir_weight[102][72],
reservoir_weight[102][73],
reservoir_weight[102][74],
reservoir_weight[102][75],
reservoir_weight[102][76],
reservoir_weight[102][77],
reservoir_weight[102][78],
reservoir_weight[102][79],
reservoir_weight[102][80],
reservoir_weight[102][81],
reservoir_weight[102][82],
reservoir_weight[102][83],
reservoir_weight[102][84],
reservoir_weight[102][85],
reservoir_weight[102][86],
reservoir_weight[102][87],
reservoir_weight[102][88],
reservoir_weight[102][89],
reservoir_weight[102][90],
reservoir_weight[102][91],
reservoir_weight[102][92],
reservoir_weight[102][93],
reservoir_weight[102][94],
reservoir_weight[102][95],
reservoir_weight[102][96],
reservoir_weight[102][97],
reservoir_weight[102][98],
reservoir_weight[102][99],
reservoir_weight[102][100],
reservoir_weight[102][101],
reservoir_weight[102][102],
reservoir_weight[102][103],
reservoir_weight[102][104],
reservoir_weight[102][105],
reservoir_weight[102][106],
reservoir_weight[102][107],
reservoir_weight[102][108],
reservoir_weight[102][109],
reservoir_weight[102][110],
reservoir_weight[102][111],
reservoir_weight[102][112],
reservoir_weight[102][113],
reservoir_weight[102][114],
reservoir_weight[102][115],
reservoir_weight[102][116],
reservoir_weight[102][117],
reservoir_weight[102][118],
reservoir_weight[102][119],
reservoir_weight[102][120],
reservoir_weight[102][121],
reservoir_weight[102][122],
reservoir_weight[102][123],
reservoir_weight[102][124],
reservoir_weight[102][125],
reservoir_weight[102][126],
reservoir_weight[102][127],
reservoir_weight[102][128],
reservoir_weight[102][129],
reservoir_weight[102][130],
reservoir_weight[102][131],
reservoir_weight[102][132],
reservoir_weight[102][133],
reservoir_weight[102][134],
reservoir_weight[102][135],
reservoir_weight[102][136],
reservoir_weight[102][137],
reservoir_weight[102][138],
reservoir_weight[102][139],
reservoir_weight[102][140],
reservoir_weight[102][141],
reservoir_weight[102][142],
reservoir_weight[102][143],
reservoir_weight[102][144],
reservoir_weight[102][145],
reservoir_weight[102][146],
reservoir_weight[102][147],
reservoir_weight[102][148],
reservoir_weight[102][149],
reservoir_weight[102][150],
reservoir_weight[102][151],
reservoir_weight[102][152],
reservoir_weight[102][153],
reservoir_weight[102][154],
reservoir_weight[102][155],
reservoir_weight[102][156],
reservoir_weight[102][157],
reservoir_weight[102][158],
reservoir_weight[102][159],
reservoir_weight[102][160],
reservoir_weight[102][161],
reservoir_weight[102][162],
reservoir_weight[102][163],
reservoir_weight[102][164],
reservoir_weight[102][165],
reservoir_weight[102][166],
reservoir_weight[102][167],
reservoir_weight[102][168],
reservoir_weight[102][169],
reservoir_weight[102][170],
reservoir_weight[102][171],
reservoir_weight[102][172],
reservoir_weight[102][173],
reservoir_weight[102][174],
reservoir_weight[102][175],
reservoir_weight[102][176],
reservoir_weight[102][177],
reservoir_weight[102][178],
reservoir_weight[102][179],
reservoir_weight[102][180],
reservoir_weight[102][181],
reservoir_weight[102][182],
reservoir_weight[102][183],
reservoir_weight[102][184],
reservoir_weight[102][185],
reservoir_weight[102][186],
reservoir_weight[102][187],
reservoir_weight[102][188],
reservoir_weight[102][189],
reservoir_weight[102][190],
reservoir_weight[102][191],
reservoir_weight[102][192],
reservoir_weight[102][193],
reservoir_weight[102][194],
reservoir_weight[102][195],
reservoir_weight[102][196],
reservoir_weight[102][197],
reservoir_weight[102][198],
reservoir_weight[102][199]
},
{reservoir_weight[103][0],
reservoir_weight[103][1],
reservoir_weight[103][2],
reservoir_weight[103][3],
reservoir_weight[103][4],
reservoir_weight[103][5],
reservoir_weight[103][6],
reservoir_weight[103][7],
reservoir_weight[103][8],
reservoir_weight[103][9],
reservoir_weight[103][10],
reservoir_weight[103][11],
reservoir_weight[103][12],
reservoir_weight[103][13],
reservoir_weight[103][14],
reservoir_weight[103][15],
reservoir_weight[103][16],
reservoir_weight[103][17],
reservoir_weight[103][18],
reservoir_weight[103][19],
reservoir_weight[103][20],
reservoir_weight[103][21],
reservoir_weight[103][22],
reservoir_weight[103][23],
reservoir_weight[103][24],
reservoir_weight[103][25],
reservoir_weight[103][26],
reservoir_weight[103][27],
reservoir_weight[103][28],
reservoir_weight[103][29],
reservoir_weight[103][30],
reservoir_weight[103][31],
reservoir_weight[103][32],
reservoir_weight[103][33],
reservoir_weight[103][34],
reservoir_weight[103][35],
reservoir_weight[103][36],
reservoir_weight[103][37],
reservoir_weight[103][38],
reservoir_weight[103][39],
reservoir_weight[103][40],
reservoir_weight[103][41],
reservoir_weight[103][42],
reservoir_weight[103][43],
reservoir_weight[103][44],
reservoir_weight[103][45],
reservoir_weight[103][46],
reservoir_weight[103][47],
reservoir_weight[103][48],
reservoir_weight[103][49],
reservoir_weight[103][50],
reservoir_weight[103][51],
reservoir_weight[103][52],
reservoir_weight[103][53],
reservoir_weight[103][54],
reservoir_weight[103][55],
reservoir_weight[103][56],
reservoir_weight[103][57],
reservoir_weight[103][58],
reservoir_weight[103][59],
reservoir_weight[103][60],
reservoir_weight[103][61],
reservoir_weight[103][62],
reservoir_weight[103][63],
reservoir_weight[103][64],
reservoir_weight[103][65],
reservoir_weight[103][66],
reservoir_weight[103][67],
reservoir_weight[103][68],
reservoir_weight[103][69],
reservoir_weight[103][70],
reservoir_weight[103][71],
reservoir_weight[103][72],
reservoir_weight[103][73],
reservoir_weight[103][74],
reservoir_weight[103][75],
reservoir_weight[103][76],
reservoir_weight[103][77],
reservoir_weight[103][78],
reservoir_weight[103][79],
reservoir_weight[103][80],
reservoir_weight[103][81],
reservoir_weight[103][82],
reservoir_weight[103][83],
reservoir_weight[103][84],
reservoir_weight[103][85],
reservoir_weight[103][86],
reservoir_weight[103][87],
reservoir_weight[103][88],
reservoir_weight[103][89],
reservoir_weight[103][90],
reservoir_weight[103][91],
reservoir_weight[103][92],
reservoir_weight[103][93],
reservoir_weight[103][94],
reservoir_weight[103][95],
reservoir_weight[103][96],
reservoir_weight[103][97],
reservoir_weight[103][98],
reservoir_weight[103][99],
reservoir_weight[103][100],
reservoir_weight[103][101],
reservoir_weight[103][102],
reservoir_weight[103][103],
reservoir_weight[103][104],
reservoir_weight[103][105],
reservoir_weight[103][106],
reservoir_weight[103][107],
reservoir_weight[103][108],
reservoir_weight[103][109],
reservoir_weight[103][110],
reservoir_weight[103][111],
reservoir_weight[103][112],
reservoir_weight[103][113],
reservoir_weight[103][114],
reservoir_weight[103][115],
reservoir_weight[103][116],
reservoir_weight[103][117],
reservoir_weight[103][118],
reservoir_weight[103][119],
reservoir_weight[103][120],
reservoir_weight[103][121],
reservoir_weight[103][122],
reservoir_weight[103][123],
reservoir_weight[103][124],
reservoir_weight[103][125],
reservoir_weight[103][126],
reservoir_weight[103][127],
reservoir_weight[103][128],
reservoir_weight[103][129],
reservoir_weight[103][130],
reservoir_weight[103][131],
reservoir_weight[103][132],
reservoir_weight[103][133],
reservoir_weight[103][134],
reservoir_weight[103][135],
reservoir_weight[103][136],
reservoir_weight[103][137],
reservoir_weight[103][138],
reservoir_weight[103][139],
reservoir_weight[103][140],
reservoir_weight[103][141],
reservoir_weight[103][142],
reservoir_weight[103][143],
reservoir_weight[103][144],
reservoir_weight[103][145],
reservoir_weight[103][146],
reservoir_weight[103][147],
reservoir_weight[103][148],
reservoir_weight[103][149],
reservoir_weight[103][150],
reservoir_weight[103][151],
reservoir_weight[103][152],
reservoir_weight[103][153],
reservoir_weight[103][154],
reservoir_weight[103][155],
reservoir_weight[103][156],
reservoir_weight[103][157],
reservoir_weight[103][158],
reservoir_weight[103][159],
reservoir_weight[103][160],
reservoir_weight[103][161],
reservoir_weight[103][162],
reservoir_weight[103][163],
reservoir_weight[103][164],
reservoir_weight[103][165],
reservoir_weight[103][166],
reservoir_weight[103][167],
reservoir_weight[103][168],
reservoir_weight[103][169],
reservoir_weight[103][170],
reservoir_weight[103][171],
reservoir_weight[103][172],
reservoir_weight[103][173],
reservoir_weight[103][174],
reservoir_weight[103][175],
reservoir_weight[103][176],
reservoir_weight[103][177],
reservoir_weight[103][178],
reservoir_weight[103][179],
reservoir_weight[103][180],
reservoir_weight[103][181],
reservoir_weight[103][182],
reservoir_weight[103][183],
reservoir_weight[103][184],
reservoir_weight[103][185],
reservoir_weight[103][186],
reservoir_weight[103][187],
reservoir_weight[103][188],
reservoir_weight[103][189],
reservoir_weight[103][190],
reservoir_weight[103][191],
reservoir_weight[103][192],
reservoir_weight[103][193],
reservoir_weight[103][194],
reservoir_weight[103][195],
reservoir_weight[103][196],
reservoir_weight[103][197],
reservoir_weight[103][198],
reservoir_weight[103][199]
},
{reservoir_weight[104][0],
reservoir_weight[104][1],
reservoir_weight[104][2],
reservoir_weight[104][3],
reservoir_weight[104][4],
reservoir_weight[104][5],
reservoir_weight[104][6],
reservoir_weight[104][7],
reservoir_weight[104][8],
reservoir_weight[104][9],
reservoir_weight[104][10],
reservoir_weight[104][11],
reservoir_weight[104][12],
reservoir_weight[104][13],
reservoir_weight[104][14],
reservoir_weight[104][15],
reservoir_weight[104][16],
reservoir_weight[104][17],
reservoir_weight[104][18],
reservoir_weight[104][19],
reservoir_weight[104][20],
reservoir_weight[104][21],
reservoir_weight[104][22],
reservoir_weight[104][23],
reservoir_weight[104][24],
reservoir_weight[104][25],
reservoir_weight[104][26],
reservoir_weight[104][27],
reservoir_weight[104][28],
reservoir_weight[104][29],
reservoir_weight[104][30],
reservoir_weight[104][31],
reservoir_weight[104][32],
reservoir_weight[104][33],
reservoir_weight[104][34],
reservoir_weight[104][35],
reservoir_weight[104][36],
reservoir_weight[104][37],
reservoir_weight[104][38],
reservoir_weight[104][39],
reservoir_weight[104][40],
reservoir_weight[104][41],
reservoir_weight[104][42],
reservoir_weight[104][43],
reservoir_weight[104][44],
reservoir_weight[104][45],
reservoir_weight[104][46],
reservoir_weight[104][47],
reservoir_weight[104][48],
reservoir_weight[104][49],
reservoir_weight[104][50],
reservoir_weight[104][51],
reservoir_weight[104][52],
reservoir_weight[104][53],
reservoir_weight[104][54],
reservoir_weight[104][55],
reservoir_weight[104][56],
reservoir_weight[104][57],
reservoir_weight[104][58],
reservoir_weight[104][59],
reservoir_weight[104][60],
reservoir_weight[104][61],
reservoir_weight[104][62],
reservoir_weight[104][63],
reservoir_weight[104][64],
reservoir_weight[104][65],
reservoir_weight[104][66],
reservoir_weight[104][67],
reservoir_weight[104][68],
reservoir_weight[104][69],
reservoir_weight[104][70],
reservoir_weight[104][71],
reservoir_weight[104][72],
reservoir_weight[104][73],
reservoir_weight[104][74],
reservoir_weight[104][75],
reservoir_weight[104][76],
reservoir_weight[104][77],
reservoir_weight[104][78],
reservoir_weight[104][79],
reservoir_weight[104][80],
reservoir_weight[104][81],
reservoir_weight[104][82],
reservoir_weight[104][83],
reservoir_weight[104][84],
reservoir_weight[104][85],
reservoir_weight[104][86],
reservoir_weight[104][87],
reservoir_weight[104][88],
reservoir_weight[104][89],
reservoir_weight[104][90],
reservoir_weight[104][91],
reservoir_weight[104][92],
reservoir_weight[104][93],
reservoir_weight[104][94],
reservoir_weight[104][95],
reservoir_weight[104][96],
reservoir_weight[104][97],
reservoir_weight[104][98],
reservoir_weight[104][99],
reservoir_weight[104][100],
reservoir_weight[104][101],
reservoir_weight[104][102],
reservoir_weight[104][103],
reservoir_weight[104][104],
reservoir_weight[104][105],
reservoir_weight[104][106],
reservoir_weight[104][107],
reservoir_weight[104][108],
reservoir_weight[104][109],
reservoir_weight[104][110],
reservoir_weight[104][111],
reservoir_weight[104][112],
reservoir_weight[104][113],
reservoir_weight[104][114],
reservoir_weight[104][115],
reservoir_weight[104][116],
reservoir_weight[104][117],
reservoir_weight[104][118],
reservoir_weight[104][119],
reservoir_weight[104][120],
reservoir_weight[104][121],
reservoir_weight[104][122],
reservoir_weight[104][123],
reservoir_weight[104][124],
reservoir_weight[104][125],
reservoir_weight[104][126],
reservoir_weight[104][127],
reservoir_weight[104][128],
reservoir_weight[104][129],
reservoir_weight[104][130],
reservoir_weight[104][131],
reservoir_weight[104][132],
reservoir_weight[104][133],
reservoir_weight[104][134],
reservoir_weight[104][135],
reservoir_weight[104][136],
reservoir_weight[104][137],
reservoir_weight[104][138],
reservoir_weight[104][139],
reservoir_weight[104][140],
reservoir_weight[104][141],
reservoir_weight[104][142],
reservoir_weight[104][143],
reservoir_weight[104][144],
reservoir_weight[104][145],
reservoir_weight[104][146],
reservoir_weight[104][147],
reservoir_weight[104][148],
reservoir_weight[104][149],
reservoir_weight[104][150],
reservoir_weight[104][151],
reservoir_weight[104][152],
reservoir_weight[104][153],
reservoir_weight[104][154],
reservoir_weight[104][155],
reservoir_weight[104][156],
reservoir_weight[104][157],
reservoir_weight[104][158],
reservoir_weight[104][159],
reservoir_weight[104][160],
reservoir_weight[104][161],
reservoir_weight[104][162],
reservoir_weight[104][163],
reservoir_weight[104][164],
reservoir_weight[104][165],
reservoir_weight[104][166],
reservoir_weight[104][167],
reservoir_weight[104][168],
reservoir_weight[104][169],
reservoir_weight[104][170],
reservoir_weight[104][171],
reservoir_weight[104][172],
reservoir_weight[104][173],
reservoir_weight[104][174],
reservoir_weight[104][175],
reservoir_weight[104][176],
reservoir_weight[104][177],
reservoir_weight[104][178],
reservoir_weight[104][179],
reservoir_weight[104][180],
reservoir_weight[104][181],
reservoir_weight[104][182],
reservoir_weight[104][183],
reservoir_weight[104][184],
reservoir_weight[104][185],
reservoir_weight[104][186],
reservoir_weight[104][187],
reservoir_weight[104][188],
reservoir_weight[104][189],
reservoir_weight[104][190],
reservoir_weight[104][191],
reservoir_weight[104][192],
reservoir_weight[104][193],
reservoir_weight[104][194],
reservoir_weight[104][195],
reservoir_weight[104][196],
reservoir_weight[104][197],
reservoir_weight[104][198],
reservoir_weight[104][199]
},
{reservoir_weight[105][0],
reservoir_weight[105][1],
reservoir_weight[105][2],
reservoir_weight[105][3],
reservoir_weight[105][4],
reservoir_weight[105][5],
reservoir_weight[105][6],
reservoir_weight[105][7],
reservoir_weight[105][8],
reservoir_weight[105][9],
reservoir_weight[105][10],
reservoir_weight[105][11],
reservoir_weight[105][12],
reservoir_weight[105][13],
reservoir_weight[105][14],
reservoir_weight[105][15],
reservoir_weight[105][16],
reservoir_weight[105][17],
reservoir_weight[105][18],
reservoir_weight[105][19],
reservoir_weight[105][20],
reservoir_weight[105][21],
reservoir_weight[105][22],
reservoir_weight[105][23],
reservoir_weight[105][24],
reservoir_weight[105][25],
reservoir_weight[105][26],
reservoir_weight[105][27],
reservoir_weight[105][28],
reservoir_weight[105][29],
reservoir_weight[105][30],
reservoir_weight[105][31],
reservoir_weight[105][32],
reservoir_weight[105][33],
reservoir_weight[105][34],
reservoir_weight[105][35],
reservoir_weight[105][36],
reservoir_weight[105][37],
reservoir_weight[105][38],
reservoir_weight[105][39],
reservoir_weight[105][40],
reservoir_weight[105][41],
reservoir_weight[105][42],
reservoir_weight[105][43],
reservoir_weight[105][44],
reservoir_weight[105][45],
reservoir_weight[105][46],
reservoir_weight[105][47],
reservoir_weight[105][48],
reservoir_weight[105][49],
reservoir_weight[105][50],
reservoir_weight[105][51],
reservoir_weight[105][52],
reservoir_weight[105][53],
reservoir_weight[105][54],
reservoir_weight[105][55],
reservoir_weight[105][56],
reservoir_weight[105][57],
reservoir_weight[105][58],
reservoir_weight[105][59],
reservoir_weight[105][60],
reservoir_weight[105][61],
reservoir_weight[105][62],
reservoir_weight[105][63],
reservoir_weight[105][64],
reservoir_weight[105][65],
reservoir_weight[105][66],
reservoir_weight[105][67],
reservoir_weight[105][68],
reservoir_weight[105][69],
reservoir_weight[105][70],
reservoir_weight[105][71],
reservoir_weight[105][72],
reservoir_weight[105][73],
reservoir_weight[105][74],
reservoir_weight[105][75],
reservoir_weight[105][76],
reservoir_weight[105][77],
reservoir_weight[105][78],
reservoir_weight[105][79],
reservoir_weight[105][80],
reservoir_weight[105][81],
reservoir_weight[105][82],
reservoir_weight[105][83],
reservoir_weight[105][84],
reservoir_weight[105][85],
reservoir_weight[105][86],
reservoir_weight[105][87],
reservoir_weight[105][88],
reservoir_weight[105][89],
reservoir_weight[105][90],
reservoir_weight[105][91],
reservoir_weight[105][92],
reservoir_weight[105][93],
reservoir_weight[105][94],
reservoir_weight[105][95],
reservoir_weight[105][96],
reservoir_weight[105][97],
reservoir_weight[105][98],
reservoir_weight[105][99],
reservoir_weight[105][100],
reservoir_weight[105][101],
reservoir_weight[105][102],
reservoir_weight[105][103],
reservoir_weight[105][104],
reservoir_weight[105][105],
reservoir_weight[105][106],
reservoir_weight[105][107],
reservoir_weight[105][108],
reservoir_weight[105][109],
reservoir_weight[105][110],
reservoir_weight[105][111],
reservoir_weight[105][112],
reservoir_weight[105][113],
reservoir_weight[105][114],
reservoir_weight[105][115],
reservoir_weight[105][116],
reservoir_weight[105][117],
reservoir_weight[105][118],
reservoir_weight[105][119],
reservoir_weight[105][120],
reservoir_weight[105][121],
reservoir_weight[105][122],
reservoir_weight[105][123],
reservoir_weight[105][124],
reservoir_weight[105][125],
reservoir_weight[105][126],
reservoir_weight[105][127],
reservoir_weight[105][128],
reservoir_weight[105][129],
reservoir_weight[105][130],
reservoir_weight[105][131],
reservoir_weight[105][132],
reservoir_weight[105][133],
reservoir_weight[105][134],
reservoir_weight[105][135],
reservoir_weight[105][136],
reservoir_weight[105][137],
reservoir_weight[105][138],
reservoir_weight[105][139],
reservoir_weight[105][140],
reservoir_weight[105][141],
reservoir_weight[105][142],
reservoir_weight[105][143],
reservoir_weight[105][144],
reservoir_weight[105][145],
reservoir_weight[105][146],
reservoir_weight[105][147],
reservoir_weight[105][148],
reservoir_weight[105][149],
reservoir_weight[105][150],
reservoir_weight[105][151],
reservoir_weight[105][152],
reservoir_weight[105][153],
reservoir_weight[105][154],
reservoir_weight[105][155],
reservoir_weight[105][156],
reservoir_weight[105][157],
reservoir_weight[105][158],
reservoir_weight[105][159],
reservoir_weight[105][160],
reservoir_weight[105][161],
reservoir_weight[105][162],
reservoir_weight[105][163],
reservoir_weight[105][164],
reservoir_weight[105][165],
reservoir_weight[105][166],
reservoir_weight[105][167],
reservoir_weight[105][168],
reservoir_weight[105][169],
reservoir_weight[105][170],
reservoir_weight[105][171],
reservoir_weight[105][172],
reservoir_weight[105][173],
reservoir_weight[105][174],
reservoir_weight[105][175],
reservoir_weight[105][176],
reservoir_weight[105][177],
reservoir_weight[105][178],
reservoir_weight[105][179],
reservoir_weight[105][180],
reservoir_weight[105][181],
reservoir_weight[105][182],
reservoir_weight[105][183],
reservoir_weight[105][184],
reservoir_weight[105][185],
reservoir_weight[105][186],
reservoir_weight[105][187],
reservoir_weight[105][188],
reservoir_weight[105][189],
reservoir_weight[105][190],
reservoir_weight[105][191],
reservoir_weight[105][192],
reservoir_weight[105][193],
reservoir_weight[105][194],
reservoir_weight[105][195],
reservoir_weight[105][196],
reservoir_weight[105][197],
reservoir_weight[105][198],
reservoir_weight[105][199]
},
{reservoir_weight[106][0],
reservoir_weight[106][1],
reservoir_weight[106][2],
reservoir_weight[106][3],
reservoir_weight[106][4],
reservoir_weight[106][5],
reservoir_weight[106][6],
reservoir_weight[106][7],
reservoir_weight[106][8],
reservoir_weight[106][9],
reservoir_weight[106][10],
reservoir_weight[106][11],
reservoir_weight[106][12],
reservoir_weight[106][13],
reservoir_weight[106][14],
reservoir_weight[106][15],
reservoir_weight[106][16],
reservoir_weight[106][17],
reservoir_weight[106][18],
reservoir_weight[106][19],
reservoir_weight[106][20],
reservoir_weight[106][21],
reservoir_weight[106][22],
reservoir_weight[106][23],
reservoir_weight[106][24],
reservoir_weight[106][25],
reservoir_weight[106][26],
reservoir_weight[106][27],
reservoir_weight[106][28],
reservoir_weight[106][29],
reservoir_weight[106][30],
reservoir_weight[106][31],
reservoir_weight[106][32],
reservoir_weight[106][33],
reservoir_weight[106][34],
reservoir_weight[106][35],
reservoir_weight[106][36],
reservoir_weight[106][37],
reservoir_weight[106][38],
reservoir_weight[106][39],
reservoir_weight[106][40],
reservoir_weight[106][41],
reservoir_weight[106][42],
reservoir_weight[106][43],
reservoir_weight[106][44],
reservoir_weight[106][45],
reservoir_weight[106][46],
reservoir_weight[106][47],
reservoir_weight[106][48],
reservoir_weight[106][49],
reservoir_weight[106][50],
reservoir_weight[106][51],
reservoir_weight[106][52],
reservoir_weight[106][53],
reservoir_weight[106][54],
reservoir_weight[106][55],
reservoir_weight[106][56],
reservoir_weight[106][57],
reservoir_weight[106][58],
reservoir_weight[106][59],
reservoir_weight[106][60],
reservoir_weight[106][61],
reservoir_weight[106][62],
reservoir_weight[106][63],
reservoir_weight[106][64],
reservoir_weight[106][65],
reservoir_weight[106][66],
reservoir_weight[106][67],
reservoir_weight[106][68],
reservoir_weight[106][69],
reservoir_weight[106][70],
reservoir_weight[106][71],
reservoir_weight[106][72],
reservoir_weight[106][73],
reservoir_weight[106][74],
reservoir_weight[106][75],
reservoir_weight[106][76],
reservoir_weight[106][77],
reservoir_weight[106][78],
reservoir_weight[106][79],
reservoir_weight[106][80],
reservoir_weight[106][81],
reservoir_weight[106][82],
reservoir_weight[106][83],
reservoir_weight[106][84],
reservoir_weight[106][85],
reservoir_weight[106][86],
reservoir_weight[106][87],
reservoir_weight[106][88],
reservoir_weight[106][89],
reservoir_weight[106][90],
reservoir_weight[106][91],
reservoir_weight[106][92],
reservoir_weight[106][93],
reservoir_weight[106][94],
reservoir_weight[106][95],
reservoir_weight[106][96],
reservoir_weight[106][97],
reservoir_weight[106][98],
reservoir_weight[106][99],
reservoir_weight[106][100],
reservoir_weight[106][101],
reservoir_weight[106][102],
reservoir_weight[106][103],
reservoir_weight[106][104],
reservoir_weight[106][105],
reservoir_weight[106][106],
reservoir_weight[106][107],
reservoir_weight[106][108],
reservoir_weight[106][109],
reservoir_weight[106][110],
reservoir_weight[106][111],
reservoir_weight[106][112],
reservoir_weight[106][113],
reservoir_weight[106][114],
reservoir_weight[106][115],
reservoir_weight[106][116],
reservoir_weight[106][117],
reservoir_weight[106][118],
reservoir_weight[106][119],
reservoir_weight[106][120],
reservoir_weight[106][121],
reservoir_weight[106][122],
reservoir_weight[106][123],
reservoir_weight[106][124],
reservoir_weight[106][125],
reservoir_weight[106][126],
reservoir_weight[106][127],
reservoir_weight[106][128],
reservoir_weight[106][129],
reservoir_weight[106][130],
reservoir_weight[106][131],
reservoir_weight[106][132],
reservoir_weight[106][133],
reservoir_weight[106][134],
reservoir_weight[106][135],
reservoir_weight[106][136],
reservoir_weight[106][137],
reservoir_weight[106][138],
reservoir_weight[106][139],
reservoir_weight[106][140],
reservoir_weight[106][141],
reservoir_weight[106][142],
reservoir_weight[106][143],
reservoir_weight[106][144],
reservoir_weight[106][145],
reservoir_weight[106][146],
reservoir_weight[106][147],
reservoir_weight[106][148],
reservoir_weight[106][149],
reservoir_weight[106][150],
reservoir_weight[106][151],
reservoir_weight[106][152],
reservoir_weight[106][153],
reservoir_weight[106][154],
reservoir_weight[106][155],
reservoir_weight[106][156],
reservoir_weight[106][157],
reservoir_weight[106][158],
reservoir_weight[106][159],
reservoir_weight[106][160],
reservoir_weight[106][161],
reservoir_weight[106][162],
reservoir_weight[106][163],
reservoir_weight[106][164],
reservoir_weight[106][165],
reservoir_weight[106][166],
reservoir_weight[106][167],
reservoir_weight[106][168],
reservoir_weight[106][169],
reservoir_weight[106][170],
reservoir_weight[106][171],
reservoir_weight[106][172],
reservoir_weight[106][173],
reservoir_weight[106][174],
reservoir_weight[106][175],
reservoir_weight[106][176],
reservoir_weight[106][177],
reservoir_weight[106][178],
reservoir_weight[106][179],
reservoir_weight[106][180],
reservoir_weight[106][181],
reservoir_weight[106][182],
reservoir_weight[106][183],
reservoir_weight[106][184],
reservoir_weight[106][185],
reservoir_weight[106][186],
reservoir_weight[106][187],
reservoir_weight[106][188],
reservoir_weight[106][189],
reservoir_weight[106][190],
reservoir_weight[106][191],
reservoir_weight[106][192],
reservoir_weight[106][193],
reservoir_weight[106][194],
reservoir_weight[106][195],
reservoir_weight[106][196],
reservoir_weight[106][197],
reservoir_weight[106][198],
reservoir_weight[106][199]
},
{reservoir_weight[107][0],
reservoir_weight[107][1],
reservoir_weight[107][2],
reservoir_weight[107][3],
reservoir_weight[107][4],
reservoir_weight[107][5],
reservoir_weight[107][6],
reservoir_weight[107][7],
reservoir_weight[107][8],
reservoir_weight[107][9],
reservoir_weight[107][10],
reservoir_weight[107][11],
reservoir_weight[107][12],
reservoir_weight[107][13],
reservoir_weight[107][14],
reservoir_weight[107][15],
reservoir_weight[107][16],
reservoir_weight[107][17],
reservoir_weight[107][18],
reservoir_weight[107][19],
reservoir_weight[107][20],
reservoir_weight[107][21],
reservoir_weight[107][22],
reservoir_weight[107][23],
reservoir_weight[107][24],
reservoir_weight[107][25],
reservoir_weight[107][26],
reservoir_weight[107][27],
reservoir_weight[107][28],
reservoir_weight[107][29],
reservoir_weight[107][30],
reservoir_weight[107][31],
reservoir_weight[107][32],
reservoir_weight[107][33],
reservoir_weight[107][34],
reservoir_weight[107][35],
reservoir_weight[107][36],
reservoir_weight[107][37],
reservoir_weight[107][38],
reservoir_weight[107][39],
reservoir_weight[107][40],
reservoir_weight[107][41],
reservoir_weight[107][42],
reservoir_weight[107][43],
reservoir_weight[107][44],
reservoir_weight[107][45],
reservoir_weight[107][46],
reservoir_weight[107][47],
reservoir_weight[107][48],
reservoir_weight[107][49],
reservoir_weight[107][50],
reservoir_weight[107][51],
reservoir_weight[107][52],
reservoir_weight[107][53],
reservoir_weight[107][54],
reservoir_weight[107][55],
reservoir_weight[107][56],
reservoir_weight[107][57],
reservoir_weight[107][58],
reservoir_weight[107][59],
reservoir_weight[107][60],
reservoir_weight[107][61],
reservoir_weight[107][62],
reservoir_weight[107][63],
reservoir_weight[107][64],
reservoir_weight[107][65],
reservoir_weight[107][66],
reservoir_weight[107][67],
reservoir_weight[107][68],
reservoir_weight[107][69],
reservoir_weight[107][70],
reservoir_weight[107][71],
reservoir_weight[107][72],
reservoir_weight[107][73],
reservoir_weight[107][74],
reservoir_weight[107][75],
reservoir_weight[107][76],
reservoir_weight[107][77],
reservoir_weight[107][78],
reservoir_weight[107][79],
reservoir_weight[107][80],
reservoir_weight[107][81],
reservoir_weight[107][82],
reservoir_weight[107][83],
reservoir_weight[107][84],
reservoir_weight[107][85],
reservoir_weight[107][86],
reservoir_weight[107][87],
reservoir_weight[107][88],
reservoir_weight[107][89],
reservoir_weight[107][90],
reservoir_weight[107][91],
reservoir_weight[107][92],
reservoir_weight[107][93],
reservoir_weight[107][94],
reservoir_weight[107][95],
reservoir_weight[107][96],
reservoir_weight[107][97],
reservoir_weight[107][98],
reservoir_weight[107][99],
reservoir_weight[107][100],
reservoir_weight[107][101],
reservoir_weight[107][102],
reservoir_weight[107][103],
reservoir_weight[107][104],
reservoir_weight[107][105],
reservoir_weight[107][106],
reservoir_weight[107][107],
reservoir_weight[107][108],
reservoir_weight[107][109],
reservoir_weight[107][110],
reservoir_weight[107][111],
reservoir_weight[107][112],
reservoir_weight[107][113],
reservoir_weight[107][114],
reservoir_weight[107][115],
reservoir_weight[107][116],
reservoir_weight[107][117],
reservoir_weight[107][118],
reservoir_weight[107][119],
reservoir_weight[107][120],
reservoir_weight[107][121],
reservoir_weight[107][122],
reservoir_weight[107][123],
reservoir_weight[107][124],
reservoir_weight[107][125],
reservoir_weight[107][126],
reservoir_weight[107][127],
reservoir_weight[107][128],
reservoir_weight[107][129],
reservoir_weight[107][130],
reservoir_weight[107][131],
reservoir_weight[107][132],
reservoir_weight[107][133],
reservoir_weight[107][134],
reservoir_weight[107][135],
reservoir_weight[107][136],
reservoir_weight[107][137],
reservoir_weight[107][138],
reservoir_weight[107][139],
reservoir_weight[107][140],
reservoir_weight[107][141],
reservoir_weight[107][142],
reservoir_weight[107][143],
reservoir_weight[107][144],
reservoir_weight[107][145],
reservoir_weight[107][146],
reservoir_weight[107][147],
reservoir_weight[107][148],
reservoir_weight[107][149],
reservoir_weight[107][150],
reservoir_weight[107][151],
reservoir_weight[107][152],
reservoir_weight[107][153],
reservoir_weight[107][154],
reservoir_weight[107][155],
reservoir_weight[107][156],
reservoir_weight[107][157],
reservoir_weight[107][158],
reservoir_weight[107][159],
reservoir_weight[107][160],
reservoir_weight[107][161],
reservoir_weight[107][162],
reservoir_weight[107][163],
reservoir_weight[107][164],
reservoir_weight[107][165],
reservoir_weight[107][166],
reservoir_weight[107][167],
reservoir_weight[107][168],
reservoir_weight[107][169],
reservoir_weight[107][170],
reservoir_weight[107][171],
reservoir_weight[107][172],
reservoir_weight[107][173],
reservoir_weight[107][174],
reservoir_weight[107][175],
reservoir_weight[107][176],
reservoir_weight[107][177],
reservoir_weight[107][178],
reservoir_weight[107][179],
reservoir_weight[107][180],
reservoir_weight[107][181],
reservoir_weight[107][182],
reservoir_weight[107][183],
reservoir_weight[107][184],
reservoir_weight[107][185],
reservoir_weight[107][186],
reservoir_weight[107][187],
reservoir_weight[107][188],
reservoir_weight[107][189],
reservoir_weight[107][190],
reservoir_weight[107][191],
reservoir_weight[107][192],
reservoir_weight[107][193],
reservoir_weight[107][194],
reservoir_weight[107][195],
reservoir_weight[107][196],
reservoir_weight[107][197],
reservoir_weight[107][198],
reservoir_weight[107][199]
},
{reservoir_weight[108][0],
reservoir_weight[108][1],
reservoir_weight[108][2],
reservoir_weight[108][3],
reservoir_weight[108][4],
reservoir_weight[108][5],
reservoir_weight[108][6],
reservoir_weight[108][7],
reservoir_weight[108][8],
reservoir_weight[108][9],
reservoir_weight[108][10],
reservoir_weight[108][11],
reservoir_weight[108][12],
reservoir_weight[108][13],
reservoir_weight[108][14],
reservoir_weight[108][15],
reservoir_weight[108][16],
reservoir_weight[108][17],
reservoir_weight[108][18],
reservoir_weight[108][19],
reservoir_weight[108][20],
reservoir_weight[108][21],
reservoir_weight[108][22],
reservoir_weight[108][23],
reservoir_weight[108][24],
reservoir_weight[108][25],
reservoir_weight[108][26],
reservoir_weight[108][27],
reservoir_weight[108][28],
reservoir_weight[108][29],
reservoir_weight[108][30],
reservoir_weight[108][31],
reservoir_weight[108][32],
reservoir_weight[108][33],
reservoir_weight[108][34],
reservoir_weight[108][35],
reservoir_weight[108][36],
reservoir_weight[108][37],
reservoir_weight[108][38],
reservoir_weight[108][39],
reservoir_weight[108][40],
reservoir_weight[108][41],
reservoir_weight[108][42],
reservoir_weight[108][43],
reservoir_weight[108][44],
reservoir_weight[108][45],
reservoir_weight[108][46],
reservoir_weight[108][47],
reservoir_weight[108][48],
reservoir_weight[108][49],
reservoir_weight[108][50],
reservoir_weight[108][51],
reservoir_weight[108][52],
reservoir_weight[108][53],
reservoir_weight[108][54],
reservoir_weight[108][55],
reservoir_weight[108][56],
reservoir_weight[108][57],
reservoir_weight[108][58],
reservoir_weight[108][59],
reservoir_weight[108][60],
reservoir_weight[108][61],
reservoir_weight[108][62],
reservoir_weight[108][63],
reservoir_weight[108][64],
reservoir_weight[108][65],
reservoir_weight[108][66],
reservoir_weight[108][67],
reservoir_weight[108][68],
reservoir_weight[108][69],
reservoir_weight[108][70],
reservoir_weight[108][71],
reservoir_weight[108][72],
reservoir_weight[108][73],
reservoir_weight[108][74],
reservoir_weight[108][75],
reservoir_weight[108][76],
reservoir_weight[108][77],
reservoir_weight[108][78],
reservoir_weight[108][79],
reservoir_weight[108][80],
reservoir_weight[108][81],
reservoir_weight[108][82],
reservoir_weight[108][83],
reservoir_weight[108][84],
reservoir_weight[108][85],
reservoir_weight[108][86],
reservoir_weight[108][87],
reservoir_weight[108][88],
reservoir_weight[108][89],
reservoir_weight[108][90],
reservoir_weight[108][91],
reservoir_weight[108][92],
reservoir_weight[108][93],
reservoir_weight[108][94],
reservoir_weight[108][95],
reservoir_weight[108][96],
reservoir_weight[108][97],
reservoir_weight[108][98],
reservoir_weight[108][99],
reservoir_weight[108][100],
reservoir_weight[108][101],
reservoir_weight[108][102],
reservoir_weight[108][103],
reservoir_weight[108][104],
reservoir_weight[108][105],
reservoir_weight[108][106],
reservoir_weight[108][107],
reservoir_weight[108][108],
reservoir_weight[108][109],
reservoir_weight[108][110],
reservoir_weight[108][111],
reservoir_weight[108][112],
reservoir_weight[108][113],
reservoir_weight[108][114],
reservoir_weight[108][115],
reservoir_weight[108][116],
reservoir_weight[108][117],
reservoir_weight[108][118],
reservoir_weight[108][119],
reservoir_weight[108][120],
reservoir_weight[108][121],
reservoir_weight[108][122],
reservoir_weight[108][123],
reservoir_weight[108][124],
reservoir_weight[108][125],
reservoir_weight[108][126],
reservoir_weight[108][127],
reservoir_weight[108][128],
reservoir_weight[108][129],
reservoir_weight[108][130],
reservoir_weight[108][131],
reservoir_weight[108][132],
reservoir_weight[108][133],
reservoir_weight[108][134],
reservoir_weight[108][135],
reservoir_weight[108][136],
reservoir_weight[108][137],
reservoir_weight[108][138],
reservoir_weight[108][139],
reservoir_weight[108][140],
reservoir_weight[108][141],
reservoir_weight[108][142],
reservoir_weight[108][143],
reservoir_weight[108][144],
reservoir_weight[108][145],
reservoir_weight[108][146],
reservoir_weight[108][147],
reservoir_weight[108][148],
reservoir_weight[108][149],
reservoir_weight[108][150],
reservoir_weight[108][151],
reservoir_weight[108][152],
reservoir_weight[108][153],
reservoir_weight[108][154],
reservoir_weight[108][155],
reservoir_weight[108][156],
reservoir_weight[108][157],
reservoir_weight[108][158],
reservoir_weight[108][159],
reservoir_weight[108][160],
reservoir_weight[108][161],
reservoir_weight[108][162],
reservoir_weight[108][163],
reservoir_weight[108][164],
reservoir_weight[108][165],
reservoir_weight[108][166],
reservoir_weight[108][167],
reservoir_weight[108][168],
reservoir_weight[108][169],
reservoir_weight[108][170],
reservoir_weight[108][171],
reservoir_weight[108][172],
reservoir_weight[108][173],
reservoir_weight[108][174],
reservoir_weight[108][175],
reservoir_weight[108][176],
reservoir_weight[108][177],
reservoir_weight[108][178],
reservoir_weight[108][179],
reservoir_weight[108][180],
reservoir_weight[108][181],
reservoir_weight[108][182],
reservoir_weight[108][183],
reservoir_weight[108][184],
reservoir_weight[108][185],
reservoir_weight[108][186],
reservoir_weight[108][187],
reservoir_weight[108][188],
reservoir_weight[108][189],
reservoir_weight[108][190],
reservoir_weight[108][191],
reservoir_weight[108][192],
reservoir_weight[108][193],
reservoir_weight[108][194],
reservoir_weight[108][195],
reservoir_weight[108][196],
reservoir_weight[108][197],
reservoir_weight[108][198],
reservoir_weight[108][199]
},
{reservoir_weight[109][0],
reservoir_weight[109][1],
reservoir_weight[109][2],
reservoir_weight[109][3],
reservoir_weight[109][4],
reservoir_weight[109][5],
reservoir_weight[109][6],
reservoir_weight[109][7],
reservoir_weight[109][8],
reservoir_weight[109][9],
reservoir_weight[109][10],
reservoir_weight[109][11],
reservoir_weight[109][12],
reservoir_weight[109][13],
reservoir_weight[109][14],
reservoir_weight[109][15],
reservoir_weight[109][16],
reservoir_weight[109][17],
reservoir_weight[109][18],
reservoir_weight[109][19],
reservoir_weight[109][20],
reservoir_weight[109][21],
reservoir_weight[109][22],
reservoir_weight[109][23],
reservoir_weight[109][24],
reservoir_weight[109][25],
reservoir_weight[109][26],
reservoir_weight[109][27],
reservoir_weight[109][28],
reservoir_weight[109][29],
reservoir_weight[109][30],
reservoir_weight[109][31],
reservoir_weight[109][32],
reservoir_weight[109][33],
reservoir_weight[109][34],
reservoir_weight[109][35],
reservoir_weight[109][36],
reservoir_weight[109][37],
reservoir_weight[109][38],
reservoir_weight[109][39],
reservoir_weight[109][40],
reservoir_weight[109][41],
reservoir_weight[109][42],
reservoir_weight[109][43],
reservoir_weight[109][44],
reservoir_weight[109][45],
reservoir_weight[109][46],
reservoir_weight[109][47],
reservoir_weight[109][48],
reservoir_weight[109][49],
reservoir_weight[109][50],
reservoir_weight[109][51],
reservoir_weight[109][52],
reservoir_weight[109][53],
reservoir_weight[109][54],
reservoir_weight[109][55],
reservoir_weight[109][56],
reservoir_weight[109][57],
reservoir_weight[109][58],
reservoir_weight[109][59],
reservoir_weight[109][60],
reservoir_weight[109][61],
reservoir_weight[109][62],
reservoir_weight[109][63],
reservoir_weight[109][64],
reservoir_weight[109][65],
reservoir_weight[109][66],
reservoir_weight[109][67],
reservoir_weight[109][68],
reservoir_weight[109][69],
reservoir_weight[109][70],
reservoir_weight[109][71],
reservoir_weight[109][72],
reservoir_weight[109][73],
reservoir_weight[109][74],
reservoir_weight[109][75],
reservoir_weight[109][76],
reservoir_weight[109][77],
reservoir_weight[109][78],
reservoir_weight[109][79],
reservoir_weight[109][80],
reservoir_weight[109][81],
reservoir_weight[109][82],
reservoir_weight[109][83],
reservoir_weight[109][84],
reservoir_weight[109][85],
reservoir_weight[109][86],
reservoir_weight[109][87],
reservoir_weight[109][88],
reservoir_weight[109][89],
reservoir_weight[109][90],
reservoir_weight[109][91],
reservoir_weight[109][92],
reservoir_weight[109][93],
reservoir_weight[109][94],
reservoir_weight[109][95],
reservoir_weight[109][96],
reservoir_weight[109][97],
reservoir_weight[109][98],
reservoir_weight[109][99],
reservoir_weight[109][100],
reservoir_weight[109][101],
reservoir_weight[109][102],
reservoir_weight[109][103],
reservoir_weight[109][104],
reservoir_weight[109][105],
reservoir_weight[109][106],
reservoir_weight[109][107],
reservoir_weight[109][108],
reservoir_weight[109][109],
reservoir_weight[109][110],
reservoir_weight[109][111],
reservoir_weight[109][112],
reservoir_weight[109][113],
reservoir_weight[109][114],
reservoir_weight[109][115],
reservoir_weight[109][116],
reservoir_weight[109][117],
reservoir_weight[109][118],
reservoir_weight[109][119],
reservoir_weight[109][120],
reservoir_weight[109][121],
reservoir_weight[109][122],
reservoir_weight[109][123],
reservoir_weight[109][124],
reservoir_weight[109][125],
reservoir_weight[109][126],
reservoir_weight[109][127],
reservoir_weight[109][128],
reservoir_weight[109][129],
reservoir_weight[109][130],
reservoir_weight[109][131],
reservoir_weight[109][132],
reservoir_weight[109][133],
reservoir_weight[109][134],
reservoir_weight[109][135],
reservoir_weight[109][136],
reservoir_weight[109][137],
reservoir_weight[109][138],
reservoir_weight[109][139],
reservoir_weight[109][140],
reservoir_weight[109][141],
reservoir_weight[109][142],
reservoir_weight[109][143],
reservoir_weight[109][144],
reservoir_weight[109][145],
reservoir_weight[109][146],
reservoir_weight[109][147],
reservoir_weight[109][148],
reservoir_weight[109][149],
reservoir_weight[109][150],
reservoir_weight[109][151],
reservoir_weight[109][152],
reservoir_weight[109][153],
reservoir_weight[109][154],
reservoir_weight[109][155],
reservoir_weight[109][156],
reservoir_weight[109][157],
reservoir_weight[109][158],
reservoir_weight[109][159],
reservoir_weight[109][160],
reservoir_weight[109][161],
reservoir_weight[109][162],
reservoir_weight[109][163],
reservoir_weight[109][164],
reservoir_weight[109][165],
reservoir_weight[109][166],
reservoir_weight[109][167],
reservoir_weight[109][168],
reservoir_weight[109][169],
reservoir_weight[109][170],
reservoir_weight[109][171],
reservoir_weight[109][172],
reservoir_weight[109][173],
reservoir_weight[109][174],
reservoir_weight[109][175],
reservoir_weight[109][176],
reservoir_weight[109][177],
reservoir_weight[109][178],
reservoir_weight[109][179],
reservoir_weight[109][180],
reservoir_weight[109][181],
reservoir_weight[109][182],
reservoir_weight[109][183],
reservoir_weight[109][184],
reservoir_weight[109][185],
reservoir_weight[109][186],
reservoir_weight[109][187],
reservoir_weight[109][188],
reservoir_weight[109][189],
reservoir_weight[109][190],
reservoir_weight[109][191],
reservoir_weight[109][192],
reservoir_weight[109][193],
reservoir_weight[109][194],
reservoir_weight[109][195],
reservoir_weight[109][196],
reservoir_weight[109][197],
reservoir_weight[109][198],
reservoir_weight[109][199]
},
{reservoir_weight[110][0],
reservoir_weight[110][1],
reservoir_weight[110][2],
reservoir_weight[110][3],
reservoir_weight[110][4],
reservoir_weight[110][5],
reservoir_weight[110][6],
reservoir_weight[110][7],
reservoir_weight[110][8],
reservoir_weight[110][9],
reservoir_weight[110][10],
reservoir_weight[110][11],
reservoir_weight[110][12],
reservoir_weight[110][13],
reservoir_weight[110][14],
reservoir_weight[110][15],
reservoir_weight[110][16],
reservoir_weight[110][17],
reservoir_weight[110][18],
reservoir_weight[110][19],
reservoir_weight[110][20],
reservoir_weight[110][21],
reservoir_weight[110][22],
reservoir_weight[110][23],
reservoir_weight[110][24],
reservoir_weight[110][25],
reservoir_weight[110][26],
reservoir_weight[110][27],
reservoir_weight[110][28],
reservoir_weight[110][29],
reservoir_weight[110][30],
reservoir_weight[110][31],
reservoir_weight[110][32],
reservoir_weight[110][33],
reservoir_weight[110][34],
reservoir_weight[110][35],
reservoir_weight[110][36],
reservoir_weight[110][37],
reservoir_weight[110][38],
reservoir_weight[110][39],
reservoir_weight[110][40],
reservoir_weight[110][41],
reservoir_weight[110][42],
reservoir_weight[110][43],
reservoir_weight[110][44],
reservoir_weight[110][45],
reservoir_weight[110][46],
reservoir_weight[110][47],
reservoir_weight[110][48],
reservoir_weight[110][49],
reservoir_weight[110][50],
reservoir_weight[110][51],
reservoir_weight[110][52],
reservoir_weight[110][53],
reservoir_weight[110][54],
reservoir_weight[110][55],
reservoir_weight[110][56],
reservoir_weight[110][57],
reservoir_weight[110][58],
reservoir_weight[110][59],
reservoir_weight[110][60],
reservoir_weight[110][61],
reservoir_weight[110][62],
reservoir_weight[110][63],
reservoir_weight[110][64],
reservoir_weight[110][65],
reservoir_weight[110][66],
reservoir_weight[110][67],
reservoir_weight[110][68],
reservoir_weight[110][69],
reservoir_weight[110][70],
reservoir_weight[110][71],
reservoir_weight[110][72],
reservoir_weight[110][73],
reservoir_weight[110][74],
reservoir_weight[110][75],
reservoir_weight[110][76],
reservoir_weight[110][77],
reservoir_weight[110][78],
reservoir_weight[110][79],
reservoir_weight[110][80],
reservoir_weight[110][81],
reservoir_weight[110][82],
reservoir_weight[110][83],
reservoir_weight[110][84],
reservoir_weight[110][85],
reservoir_weight[110][86],
reservoir_weight[110][87],
reservoir_weight[110][88],
reservoir_weight[110][89],
reservoir_weight[110][90],
reservoir_weight[110][91],
reservoir_weight[110][92],
reservoir_weight[110][93],
reservoir_weight[110][94],
reservoir_weight[110][95],
reservoir_weight[110][96],
reservoir_weight[110][97],
reservoir_weight[110][98],
reservoir_weight[110][99],
reservoir_weight[110][100],
reservoir_weight[110][101],
reservoir_weight[110][102],
reservoir_weight[110][103],
reservoir_weight[110][104],
reservoir_weight[110][105],
reservoir_weight[110][106],
reservoir_weight[110][107],
reservoir_weight[110][108],
reservoir_weight[110][109],
reservoir_weight[110][110],
reservoir_weight[110][111],
reservoir_weight[110][112],
reservoir_weight[110][113],
reservoir_weight[110][114],
reservoir_weight[110][115],
reservoir_weight[110][116],
reservoir_weight[110][117],
reservoir_weight[110][118],
reservoir_weight[110][119],
reservoir_weight[110][120],
reservoir_weight[110][121],
reservoir_weight[110][122],
reservoir_weight[110][123],
reservoir_weight[110][124],
reservoir_weight[110][125],
reservoir_weight[110][126],
reservoir_weight[110][127],
reservoir_weight[110][128],
reservoir_weight[110][129],
reservoir_weight[110][130],
reservoir_weight[110][131],
reservoir_weight[110][132],
reservoir_weight[110][133],
reservoir_weight[110][134],
reservoir_weight[110][135],
reservoir_weight[110][136],
reservoir_weight[110][137],
reservoir_weight[110][138],
reservoir_weight[110][139],
reservoir_weight[110][140],
reservoir_weight[110][141],
reservoir_weight[110][142],
reservoir_weight[110][143],
reservoir_weight[110][144],
reservoir_weight[110][145],
reservoir_weight[110][146],
reservoir_weight[110][147],
reservoir_weight[110][148],
reservoir_weight[110][149],
reservoir_weight[110][150],
reservoir_weight[110][151],
reservoir_weight[110][152],
reservoir_weight[110][153],
reservoir_weight[110][154],
reservoir_weight[110][155],
reservoir_weight[110][156],
reservoir_weight[110][157],
reservoir_weight[110][158],
reservoir_weight[110][159],
reservoir_weight[110][160],
reservoir_weight[110][161],
reservoir_weight[110][162],
reservoir_weight[110][163],
reservoir_weight[110][164],
reservoir_weight[110][165],
reservoir_weight[110][166],
reservoir_weight[110][167],
reservoir_weight[110][168],
reservoir_weight[110][169],
reservoir_weight[110][170],
reservoir_weight[110][171],
reservoir_weight[110][172],
reservoir_weight[110][173],
reservoir_weight[110][174],
reservoir_weight[110][175],
reservoir_weight[110][176],
reservoir_weight[110][177],
reservoir_weight[110][178],
reservoir_weight[110][179],
reservoir_weight[110][180],
reservoir_weight[110][181],
reservoir_weight[110][182],
reservoir_weight[110][183],
reservoir_weight[110][184],
reservoir_weight[110][185],
reservoir_weight[110][186],
reservoir_weight[110][187],
reservoir_weight[110][188],
reservoir_weight[110][189],
reservoir_weight[110][190],
reservoir_weight[110][191],
reservoir_weight[110][192],
reservoir_weight[110][193],
reservoir_weight[110][194],
reservoir_weight[110][195],
reservoir_weight[110][196],
reservoir_weight[110][197],
reservoir_weight[110][198],
reservoir_weight[110][199]
},
{reservoir_weight[111][0],
reservoir_weight[111][1],
reservoir_weight[111][2],
reservoir_weight[111][3],
reservoir_weight[111][4],
reservoir_weight[111][5],
reservoir_weight[111][6],
reservoir_weight[111][7],
reservoir_weight[111][8],
reservoir_weight[111][9],
reservoir_weight[111][10],
reservoir_weight[111][11],
reservoir_weight[111][12],
reservoir_weight[111][13],
reservoir_weight[111][14],
reservoir_weight[111][15],
reservoir_weight[111][16],
reservoir_weight[111][17],
reservoir_weight[111][18],
reservoir_weight[111][19],
reservoir_weight[111][20],
reservoir_weight[111][21],
reservoir_weight[111][22],
reservoir_weight[111][23],
reservoir_weight[111][24],
reservoir_weight[111][25],
reservoir_weight[111][26],
reservoir_weight[111][27],
reservoir_weight[111][28],
reservoir_weight[111][29],
reservoir_weight[111][30],
reservoir_weight[111][31],
reservoir_weight[111][32],
reservoir_weight[111][33],
reservoir_weight[111][34],
reservoir_weight[111][35],
reservoir_weight[111][36],
reservoir_weight[111][37],
reservoir_weight[111][38],
reservoir_weight[111][39],
reservoir_weight[111][40],
reservoir_weight[111][41],
reservoir_weight[111][42],
reservoir_weight[111][43],
reservoir_weight[111][44],
reservoir_weight[111][45],
reservoir_weight[111][46],
reservoir_weight[111][47],
reservoir_weight[111][48],
reservoir_weight[111][49],
reservoir_weight[111][50],
reservoir_weight[111][51],
reservoir_weight[111][52],
reservoir_weight[111][53],
reservoir_weight[111][54],
reservoir_weight[111][55],
reservoir_weight[111][56],
reservoir_weight[111][57],
reservoir_weight[111][58],
reservoir_weight[111][59],
reservoir_weight[111][60],
reservoir_weight[111][61],
reservoir_weight[111][62],
reservoir_weight[111][63],
reservoir_weight[111][64],
reservoir_weight[111][65],
reservoir_weight[111][66],
reservoir_weight[111][67],
reservoir_weight[111][68],
reservoir_weight[111][69],
reservoir_weight[111][70],
reservoir_weight[111][71],
reservoir_weight[111][72],
reservoir_weight[111][73],
reservoir_weight[111][74],
reservoir_weight[111][75],
reservoir_weight[111][76],
reservoir_weight[111][77],
reservoir_weight[111][78],
reservoir_weight[111][79],
reservoir_weight[111][80],
reservoir_weight[111][81],
reservoir_weight[111][82],
reservoir_weight[111][83],
reservoir_weight[111][84],
reservoir_weight[111][85],
reservoir_weight[111][86],
reservoir_weight[111][87],
reservoir_weight[111][88],
reservoir_weight[111][89],
reservoir_weight[111][90],
reservoir_weight[111][91],
reservoir_weight[111][92],
reservoir_weight[111][93],
reservoir_weight[111][94],
reservoir_weight[111][95],
reservoir_weight[111][96],
reservoir_weight[111][97],
reservoir_weight[111][98],
reservoir_weight[111][99],
reservoir_weight[111][100],
reservoir_weight[111][101],
reservoir_weight[111][102],
reservoir_weight[111][103],
reservoir_weight[111][104],
reservoir_weight[111][105],
reservoir_weight[111][106],
reservoir_weight[111][107],
reservoir_weight[111][108],
reservoir_weight[111][109],
reservoir_weight[111][110],
reservoir_weight[111][111],
reservoir_weight[111][112],
reservoir_weight[111][113],
reservoir_weight[111][114],
reservoir_weight[111][115],
reservoir_weight[111][116],
reservoir_weight[111][117],
reservoir_weight[111][118],
reservoir_weight[111][119],
reservoir_weight[111][120],
reservoir_weight[111][121],
reservoir_weight[111][122],
reservoir_weight[111][123],
reservoir_weight[111][124],
reservoir_weight[111][125],
reservoir_weight[111][126],
reservoir_weight[111][127],
reservoir_weight[111][128],
reservoir_weight[111][129],
reservoir_weight[111][130],
reservoir_weight[111][131],
reservoir_weight[111][132],
reservoir_weight[111][133],
reservoir_weight[111][134],
reservoir_weight[111][135],
reservoir_weight[111][136],
reservoir_weight[111][137],
reservoir_weight[111][138],
reservoir_weight[111][139],
reservoir_weight[111][140],
reservoir_weight[111][141],
reservoir_weight[111][142],
reservoir_weight[111][143],
reservoir_weight[111][144],
reservoir_weight[111][145],
reservoir_weight[111][146],
reservoir_weight[111][147],
reservoir_weight[111][148],
reservoir_weight[111][149],
reservoir_weight[111][150],
reservoir_weight[111][151],
reservoir_weight[111][152],
reservoir_weight[111][153],
reservoir_weight[111][154],
reservoir_weight[111][155],
reservoir_weight[111][156],
reservoir_weight[111][157],
reservoir_weight[111][158],
reservoir_weight[111][159],
reservoir_weight[111][160],
reservoir_weight[111][161],
reservoir_weight[111][162],
reservoir_weight[111][163],
reservoir_weight[111][164],
reservoir_weight[111][165],
reservoir_weight[111][166],
reservoir_weight[111][167],
reservoir_weight[111][168],
reservoir_weight[111][169],
reservoir_weight[111][170],
reservoir_weight[111][171],
reservoir_weight[111][172],
reservoir_weight[111][173],
reservoir_weight[111][174],
reservoir_weight[111][175],
reservoir_weight[111][176],
reservoir_weight[111][177],
reservoir_weight[111][178],
reservoir_weight[111][179],
reservoir_weight[111][180],
reservoir_weight[111][181],
reservoir_weight[111][182],
reservoir_weight[111][183],
reservoir_weight[111][184],
reservoir_weight[111][185],
reservoir_weight[111][186],
reservoir_weight[111][187],
reservoir_weight[111][188],
reservoir_weight[111][189],
reservoir_weight[111][190],
reservoir_weight[111][191],
reservoir_weight[111][192],
reservoir_weight[111][193],
reservoir_weight[111][194],
reservoir_weight[111][195],
reservoir_weight[111][196],
reservoir_weight[111][197],
reservoir_weight[111][198],
reservoir_weight[111][199]
},
{reservoir_weight[112][0],
reservoir_weight[112][1],
reservoir_weight[112][2],
reservoir_weight[112][3],
reservoir_weight[112][4],
reservoir_weight[112][5],
reservoir_weight[112][6],
reservoir_weight[112][7],
reservoir_weight[112][8],
reservoir_weight[112][9],
reservoir_weight[112][10],
reservoir_weight[112][11],
reservoir_weight[112][12],
reservoir_weight[112][13],
reservoir_weight[112][14],
reservoir_weight[112][15],
reservoir_weight[112][16],
reservoir_weight[112][17],
reservoir_weight[112][18],
reservoir_weight[112][19],
reservoir_weight[112][20],
reservoir_weight[112][21],
reservoir_weight[112][22],
reservoir_weight[112][23],
reservoir_weight[112][24],
reservoir_weight[112][25],
reservoir_weight[112][26],
reservoir_weight[112][27],
reservoir_weight[112][28],
reservoir_weight[112][29],
reservoir_weight[112][30],
reservoir_weight[112][31],
reservoir_weight[112][32],
reservoir_weight[112][33],
reservoir_weight[112][34],
reservoir_weight[112][35],
reservoir_weight[112][36],
reservoir_weight[112][37],
reservoir_weight[112][38],
reservoir_weight[112][39],
reservoir_weight[112][40],
reservoir_weight[112][41],
reservoir_weight[112][42],
reservoir_weight[112][43],
reservoir_weight[112][44],
reservoir_weight[112][45],
reservoir_weight[112][46],
reservoir_weight[112][47],
reservoir_weight[112][48],
reservoir_weight[112][49],
reservoir_weight[112][50],
reservoir_weight[112][51],
reservoir_weight[112][52],
reservoir_weight[112][53],
reservoir_weight[112][54],
reservoir_weight[112][55],
reservoir_weight[112][56],
reservoir_weight[112][57],
reservoir_weight[112][58],
reservoir_weight[112][59],
reservoir_weight[112][60],
reservoir_weight[112][61],
reservoir_weight[112][62],
reservoir_weight[112][63],
reservoir_weight[112][64],
reservoir_weight[112][65],
reservoir_weight[112][66],
reservoir_weight[112][67],
reservoir_weight[112][68],
reservoir_weight[112][69],
reservoir_weight[112][70],
reservoir_weight[112][71],
reservoir_weight[112][72],
reservoir_weight[112][73],
reservoir_weight[112][74],
reservoir_weight[112][75],
reservoir_weight[112][76],
reservoir_weight[112][77],
reservoir_weight[112][78],
reservoir_weight[112][79],
reservoir_weight[112][80],
reservoir_weight[112][81],
reservoir_weight[112][82],
reservoir_weight[112][83],
reservoir_weight[112][84],
reservoir_weight[112][85],
reservoir_weight[112][86],
reservoir_weight[112][87],
reservoir_weight[112][88],
reservoir_weight[112][89],
reservoir_weight[112][90],
reservoir_weight[112][91],
reservoir_weight[112][92],
reservoir_weight[112][93],
reservoir_weight[112][94],
reservoir_weight[112][95],
reservoir_weight[112][96],
reservoir_weight[112][97],
reservoir_weight[112][98],
reservoir_weight[112][99],
reservoir_weight[112][100],
reservoir_weight[112][101],
reservoir_weight[112][102],
reservoir_weight[112][103],
reservoir_weight[112][104],
reservoir_weight[112][105],
reservoir_weight[112][106],
reservoir_weight[112][107],
reservoir_weight[112][108],
reservoir_weight[112][109],
reservoir_weight[112][110],
reservoir_weight[112][111],
reservoir_weight[112][112],
reservoir_weight[112][113],
reservoir_weight[112][114],
reservoir_weight[112][115],
reservoir_weight[112][116],
reservoir_weight[112][117],
reservoir_weight[112][118],
reservoir_weight[112][119],
reservoir_weight[112][120],
reservoir_weight[112][121],
reservoir_weight[112][122],
reservoir_weight[112][123],
reservoir_weight[112][124],
reservoir_weight[112][125],
reservoir_weight[112][126],
reservoir_weight[112][127],
reservoir_weight[112][128],
reservoir_weight[112][129],
reservoir_weight[112][130],
reservoir_weight[112][131],
reservoir_weight[112][132],
reservoir_weight[112][133],
reservoir_weight[112][134],
reservoir_weight[112][135],
reservoir_weight[112][136],
reservoir_weight[112][137],
reservoir_weight[112][138],
reservoir_weight[112][139],
reservoir_weight[112][140],
reservoir_weight[112][141],
reservoir_weight[112][142],
reservoir_weight[112][143],
reservoir_weight[112][144],
reservoir_weight[112][145],
reservoir_weight[112][146],
reservoir_weight[112][147],
reservoir_weight[112][148],
reservoir_weight[112][149],
reservoir_weight[112][150],
reservoir_weight[112][151],
reservoir_weight[112][152],
reservoir_weight[112][153],
reservoir_weight[112][154],
reservoir_weight[112][155],
reservoir_weight[112][156],
reservoir_weight[112][157],
reservoir_weight[112][158],
reservoir_weight[112][159],
reservoir_weight[112][160],
reservoir_weight[112][161],
reservoir_weight[112][162],
reservoir_weight[112][163],
reservoir_weight[112][164],
reservoir_weight[112][165],
reservoir_weight[112][166],
reservoir_weight[112][167],
reservoir_weight[112][168],
reservoir_weight[112][169],
reservoir_weight[112][170],
reservoir_weight[112][171],
reservoir_weight[112][172],
reservoir_weight[112][173],
reservoir_weight[112][174],
reservoir_weight[112][175],
reservoir_weight[112][176],
reservoir_weight[112][177],
reservoir_weight[112][178],
reservoir_weight[112][179],
reservoir_weight[112][180],
reservoir_weight[112][181],
reservoir_weight[112][182],
reservoir_weight[112][183],
reservoir_weight[112][184],
reservoir_weight[112][185],
reservoir_weight[112][186],
reservoir_weight[112][187],
reservoir_weight[112][188],
reservoir_weight[112][189],
reservoir_weight[112][190],
reservoir_weight[112][191],
reservoir_weight[112][192],
reservoir_weight[112][193],
reservoir_weight[112][194],
reservoir_weight[112][195],
reservoir_weight[112][196],
reservoir_weight[112][197],
reservoir_weight[112][198],
reservoir_weight[112][199]
},
{reservoir_weight[113][0],
reservoir_weight[113][1],
reservoir_weight[113][2],
reservoir_weight[113][3],
reservoir_weight[113][4],
reservoir_weight[113][5],
reservoir_weight[113][6],
reservoir_weight[113][7],
reservoir_weight[113][8],
reservoir_weight[113][9],
reservoir_weight[113][10],
reservoir_weight[113][11],
reservoir_weight[113][12],
reservoir_weight[113][13],
reservoir_weight[113][14],
reservoir_weight[113][15],
reservoir_weight[113][16],
reservoir_weight[113][17],
reservoir_weight[113][18],
reservoir_weight[113][19],
reservoir_weight[113][20],
reservoir_weight[113][21],
reservoir_weight[113][22],
reservoir_weight[113][23],
reservoir_weight[113][24],
reservoir_weight[113][25],
reservoir_weight[113][26],
reservoir_weight[113][27],
reservoir_weight[113][28],
reservoir_weight[113][29],
reservoir_weight[113][30],
reservoir_weight[113][31],
reservoir_weight[113][32],
reservoir_weight[113][33],
reservoir_weight[113][34],
reservoir_weight[113][35],
reservoir_weight[113][36],
reservoir_weight[113][37],
reservoir_weight[113][38],
reservoir_weight[113][39],
reservoir_weight[113][40],
reservoir_weight[113][41],
reservoir_weight[113][42],
reservoir_weight[113][43],
reservoir_weight[113][44],
reservoir_weight[113][45],
reservoir_weight[113][46],
reservoir_weight[113][47],
reservoir_weight[113][48],
reservoir_weight[113][49],
reservoir_weight[113][50],
reservoir_weight[113][51],
reservoir_weight[113][52],
reservoir_weight[113][53],
reservoir_weight[113][54],
reservoir_weight[113][55],
reservoir_weight[113][56],
reservoir_weight[113][57],
reservoir_weight[113][58],
reservoir_weight[113][59],
reservoir_weight[113][60],
reservoir_weight[113][61],
reservoir_weight[113][62],
reservoir_weight[113][63],
reservoir_weight[113][64],
reservoir_weight[113][65],
reservoir_weight[113][66],
reservoir_weight[113][67],
reservoir_weight[113][68],
reservoir_weight[113][69],
reservoir_weight[113][70],
reservoir_weight[113][71],
reservoir_weight[113][72],
reservoir_weight[113][73],
reservoir_weight[113][74],
reservoir_weight[113][75],
reservoir_weight[113][76],
reservoir_weight[113][77],
reservoir_weight[113][78],
reservoir_weight[113][79],
reservoir_weight[113][80],
reservoir_weight[113][81],
reservoir_weight[113][82],
reservoir_weight[113][83],
reservoir_weight[113][84],
reservoir_weight[113][85],
reservoir_weight[113][86],
reservoir_weight[113][87],
reservoir_weight[113][88],
reservoir_weight[113][89],
reservoir_weight[113][90],
reservoir_weight[113][91],
reservoir_weight[113][92],
reservoir_weight[113][93],
reservoir_weight[113][94],
reservoir_weight[113][95],
reservoir_weight[113][96],
reservoir_weight[113][97],
reservoir_weight[113][98],
reservoir_weight[113][99],
reservoir_weight[113][100],
reservoir_weight[113][101],
reservoir_weight[113][102],
reservoir_weight[113][103],
reservoir_weight[113][104],
reservoir_weight[113][105],
reservoir_weight[113][106],
reservoir_weight[113][107],
reservoir_weight[113][108],
reservoir_weight[113][109],
reservoir_weight[113][110],
reservoir_weight[113][111],
reservoir_weight[113][112],
reservoir_weight[113][113],
reservoir_weight[113][114],
reservoir_weight[113][115],
reservoir_weight[113][116],
reservoir_weight[113][117],
reservoir_weight[113][118],
reservoir_weight[113][119],
reservoir_weight[113][120],
reservoir_weight[113][121],
reservoir_weight[113][122],
reservoir_weight[113][123],
reservoir_weight[113][124],
reservoir_weight[113][125],
reservoir_weight[113][126],
reservoir_weight[113][127],
reservoir_weight[113][128],
reservoir_weight[113][129],
reservoir_weight[113][130],
reservoir_weight[113][131],
reservoir_weight[113][132],
reservoir_weight[113][133],
reservoir_weight[113][134],
reservoir_weight[113][135],
reservoir_weight[113][136],
reservoir_weight[113][137],
reservoir_weight[113][138],
reservoir_weight[113][139],
reservoir_weight[113][140],
reservoir_weight[113][141],
reservoir_weight[113][142],
reservoir_weight[113][143],
reservoir_weight[113][144],
reservoir_weight[113][145],
reservoir_weight[113][146],
reservoir_weight[113][147],
reservoir_weight[113][148],
reservoir_weight[113][149],
reservoir_weight[113][150],
reservoir_weight[113][151],
reservoir_weight[113][152],
reservoir_weight[113][153],
reservoir_weight[113][154],
reservoir_weight[113][155],
reservoir_weight[113][156],
reservoir_weight[113][157],
reservoir_weight[113][158],
reservoir_weight[113][159],
reservoir_weight[113][160],
reservoir_weight[113][161],
reservoir_weight[113][162],
reservoir_weight[113][163],
reservoir_weight[113][164],
reservoir_weight[113][165],
reservoir_weight[113][166],
reservoir_weight[113][167],
reservoir_weight[113][168],
reservoir_weight[113][169],
reservoir_weight[113][170],
reservoir_weight[113][171],
reservoir_weight[113][172],
reservoir_weight[113][173],
reservoir_weight[113][174],
reservoir_weight[113][175],
reservoir_weight[113][176],
reservoir_weight[113][177],
reservoir_weight[113][178],
reservoir_weight[113][179],
reservoir_weight[113][180],
reservoir_weight[113][181],
reservoir_weight[113][182],
reservoir_weight[113][183],
reservoir_weight[113][184],
reservoir_weight[113][185],
reservoir_weight[113][186],
reservoir_weight[113][187],
reservoir_weight[113][188],
reservoir_weight[113][189],
reservoir_weight[113][190],
reservoir_weight[113][191],
reservoir_weight[113][192],
reservoir_weight[113][193],
reservoir_weight[113][194],
reservoir_weight[113][195],
reservoir_weight[113][196],
reservoir_weight[113][197],
reservoir_weight[113][198],
reservoir_weight[113][199]
},
{reservoir_weight[114][0],
reservoir_weight[114][1],
reservoir_weight[114][2],
reservoir_weight[114][3],
reservoir_weight[114][4],
reservoir_weight[114][5],
reservoir_weight[114][6],
reservoir_weight[114][7],
reservoir_weight[114][8],
reservoir_weight[114][9],
reservoir_weight[114][10],
reservoir_weight[114][11],
reservoir_weight[114][12],
reservoir_weight[114][13],
reservoir_weight[114][14],
reservoir_weight[114][15],
reservoir_weight[114][16],
reservoir_weight[114][17],
reservoir_weight[114][18],
reservoir_weight[114][19],
reservoir_weight[114][20],
reservoir_weight[114][21],
reservoir_weight[114][22],
reservoir_weight[114][23],
reservoir_weight[114][24],
reservoir_weight[114][25],
reservoir_weight[114][26],
reservoir_weight[114][27],
reservoir_weight[114][28],
reservoir_weight[114][29],
reservoir_weight[114][30],
reservoir_weight[114][31],
reservoir_weight[114][32],
reservoir_weight[114][33],
reservoir_weight[114][34],
reservoir_weight[114][35],
reservoir_weight[114][36],
reservoir_weight[114][37],
reservoir_weight[114][38],
reservoir_weight[114][39],
reservoir_weight[114][40],
reservoir_weight[114][41],
reservoir_weight[114][42],
reservoir_weight[114][43],
reservoir_weight[114][44],
reservoir_weight[114][45],
reservoir_weight[114][46],
reservoir_weight[114][47],
reservoir_weight[114][48],
reservoir_weight[114][49],
reservoir_weight[114][50],
reservoir_weight[114][51],
reservoir_weight[114][52],
reservoir_weight[114][53],
reservoir_weight[114][54],
reservoir_weight[114][55],
reservoir_weight[114][56],
reservoir_weight[114][57],
reservoir_weight[114][58],
reservoir_weight[114][59],
reservoir_weight[114][60],
reservoir_weight[114][61],
reservoir_weight[114][62],
reservoir_weight[114][63],
reservoir_weight[114][64],
reservoir_weight[114][65],
reservoir_weight[114][66],
reservoir_weight[114][67],
reservoir_weight[114][68],
reservoir_weight[114][69],
reservoir_weight[114][70],
reservoir_weight[114][71],
reservoir_weight[114][72],
reservoir_weight[114][73],
reservoir_weight[114][74],
reservoir_weight[114][75],
reservoir_weight[114][76],
reservoir_weight[114][77],
reservoir_weight[114][78],
reservoir_weight[114][79],
reservoir_weight[114][80],
reservoir_weight[114][81],
reservoir_weight[114][82],
reservoir_weight[114][83],
reservoir_weight[114][84],
reservoir_weight[114][85],
reservoir_weight[114][86],
reservoir_weight[114][87],
reservoir_weight[114][88],
reservoir_weight[114][89],
reservoir_weight[114][90],
reservoir_weight[114][91],
reservoir_weight[114][92],
reservoir_weight[114][93],
reservoir_weight[114][94],
reservoir_weight[114][95],
reservoir_weight[114][96],
reservoir_weight[114][97],
reservoir_weight[114][98],
reservoir_weight[114][99],
reservoir_weight[114][100],
reservoir_weight[114][101],
reservoir_weight[114][102],
reservoir_weight[114][103],
reservoir_weight[114][104],
reservoir_weight[114][105],
reservoir_weight[114][106],
reservoir_weight[114][107],
reservoir_weight[114][108],
reservoir_weight[114][109],
reservoir_weight[114][110],
reservoir_weight[114][111],
reservoir_weight[114][112],
reservoir_weight[114][113],
reservoir_weight[114][114],
reservoir_weight[114][115],
reservoir_weight[114][116],
reservoir_weight[114][117],
reservoir_weight[114][118],
reservoir_weight[114][119],
reservoir_weight[114][120],
reservoir_weight[114][121],
reservoir_weight[114][122],
reservoir_weight[114][123],
reservoir_weight[114][124],
reservoir_weight[114][125],
reservoir_weight[114][126],
reservoir_weight[114][127],
reservoir_weight[114][128],
reservoir_weight[114][129],
reservoir_weight[114][130],
reservoir_weight[114][131],
reservoir_weight[114][132],
reservoir_weight[114][133],
reservoir_weight[114][134],
reservoir_weight[114][135],
reservoir_weight[114][136],
reservoir_weight[114][137],
reservoir_weight[114][138],
reservoir_weight[114][139],
reservoir_weight[114][140],
reservoir_weight[114][141],
reservoir_weight[114][142],
reservoir_weight[114][143],
reservoir_weight[114][144],
reservoir_weight[114][145],
reservoir_weight[114][146],
reservoir_weight[114][147],
reservoir_weight[114][148],
reservoir_weight[114][149],
reservoir_weight[114][150],
reservoir_weight[114][151],
reservoir_weight[114][152],
reservoir_weight[114][153],
reservoir_weight[114][154],
reservoir_weight[114][155],
reservoir_weight[114][156],
reservoir_weight[114][157],
reservoir_weight[114][158],
reservoir_weight[114][159],
reservoir_weight[114][160],
reservoir_weight[114][161],
reservoir_weight[114][162],
reservoir_weight[114][163],
reservoir_weight[114][164],
reservoir_weight[114][165],
reservoir_weight[114][166],
reservoir_weight[114][167],
reservoir_weight[114][168],
reservoir_weight[114][169],
reservoir_weight[114][170],
reservoir_weight[114][171],
reservoir_weight[114][172],
reservoir_weight[114][173],
reservoir_weight[114][174],
reservoir_weight[114][175],
reservoir_weight[114][176],
reservoir_weight[114][177],
reservoir_weight[114][178],
reservoir_weight[114][179],
reservoir_weight[114][180],
reservoir_weight[114][181],
reservoir_weight[114][182],
reservoir_weight[114][183],
reservoir_weight[114][184],
reservoir_weight[114][185],
reservoir_weight[114][186],
reservoir_weight[114][187],
reservoir_weight[114][188],
reservoir_weight[114][189],
reservoir_weight[114][190],
reservoir_weight[114][191],
reservoir_weight[114][192],
reservoir_weight[114][193],
reservoir_weight[114][194],
reservoir_weight[114][195],
reservoir_weight[114][196],
reservoir_weight[114][197],
reservoir_weight[114][198],
reservoir_weight[114][199]
},
{reservoir_weight[115][0],
reservoir_weight[115][1],
reservoir_weight[115][2],
reservoir_weight[115][3],
reservoir_weight[115][4],
reservoir_weight[115][5],
reservoir_weight[115][6],
reservoir_weight[115][7],
reservoir_weight[115][8],
reservoir_weight[115][9],
reservoir_weight[115][10],
reservoir_weight[115][11],
reservoir_weight[115][12],
reservoir_weight[115][13],
reservoir_weight[115][14],
reservoir_weight[115][15],
reservoir_weight[115][16],
reservoir_weight[115][17],
reservoir_weight[115][18],
reservoir_weight[115][19],
reservoir_weight[115][20],
reservoir_weight[115][21],
reservoir_weight[115][22],
reservoir_weight[115][23],
reservoir_weight[115][24],
reservoir_weight[115][25],
reservoir_weight[115][26],
reservoir_weight[115][27],
reservoir_weight[115][28],
reservoir_weight[115][29],
reservoir_weight[115][30],
reservoir_weight[115][31],
reservoir_weight[115][32],
reservoir_weight[115][33],
reservoir_weight[115][34],
reservoir_weight[115][35],
reservoir_weight[115][36],
reservoir_weight[115][37],
reservoir_weight[115][38],
reservoir_weight[115][39],
reservoir_weight[115][40],
reservoir_weight[115][41],
reservoir_weight[115][42],
reservoir_weight[115][43],
reservoir_weight[115][44],
reservoir_weight[115][45],
reservoir_weight[115][46],
reservoir_weight[115][47],
reservoir_weight[115][48],
reservoir_weight[115][49],
reservoir_weight[115][50],
reservoir_weight[115][51],
reservoir_weight[115][52],
reservoir_weight[115][53],
reservoir_weight[115][54],
reservoir_weight[115][55],
reservoir_weight[115][56],
reservoir_weight[115][57],
reservoir_weight[115][58],
reservoir_weight[115][59],
reservoir_weight[115][60],
reservoir_weight[115][61],
reservoir_weight[115][62],
reservoir_weight[115][63],
reservoir_weight[115][64],
reservoir_weight[115][65],
reservoir_weight[115][66],
reservoir_weight[115][67],
reservoir_weight[115][68],
reservoir_weight[115][69],
reservoir_weight[115][70],
reservoir_weight[115][71],
reservoir_weight[115][72],
reservoir_weight[115][73],
reservoir_weight[115][74],
reservoir_weight[115][75],
reservoir_weight[115][76],
reservoir_weight[115][77],
reservoir_weight[115][78],
reservoir_weight[115][79],
reservoir_weight[115][80],
reservoir_weight[115][81],
reservoir_weight[115][82],
reservoir_weight[115][83],
reservoir_weight[115][84],
reservoir_weight[115][85],
reservoir_weight[115][86],
reservoir_weight[115][87],
reservoir_weight[115][88],
reservoir_weight[115][89],
reservoir_weight[115][90],
reservoir_weight[115][91],
reservoir_weight[115][92],
reservoir_weight[115][93],
reservoir_weight[115][94],
reservoir_weight[115][95],
reservoir_weight[115][96],
reservoir_weight[115][97],
reservoir_weight[115][98],
reservoir_weight[115][99],
reservoir_weight[115][100],
reservoir_weight[115][101],
reservoir_weight[115][102],
reservoir_weight[115][103],
reservoir_weight[115][104],
reservoir_weight[115][105],
reservoir_weight[115][106],
reservoir_weight[115][107],
reservoir_weight[115][108],
reservoir_weight[115][109],
reservoir_weight[115][110],
reservoir_weight[115][111],
reservoir_weight[115][112],
reservoir_weight[115][113],
reservoir_weight[115][114],
reservoir_weight[115][115],
reservoir_weight[115][116],
reservoir_weight[115][117],
reservoir_weight[115][118],
reservoir_weight[115][119],
reservoir_weight[115][120],
reservoir_weight[115][121],
reservoir_weight[115][122],
reservoir_weight[115][123],
reservoir_weight[115][124],
reservoir_weight[115][125],
reservoir_weight[115][126],
reservoir_weight[115][127],
reservoir_weight[115][128],
reservoir_weight[115][129],
reservoir_weight[115][130],
reservoir_weight[115][131],
reservoir_weight[115][132],
reservoir_weight[115][133],
reservoir_weight[115][134],
reservoir_weight[115][135],
reservoir_weight[115][136],
reservoir_weight[115][137],
reservoir_weight[115][138],
reservoir_weight[115][139],
reservoir_weight[115][140],
reservoir_weight[115][141],
reservoir_weight[115][142],
reservoir_weight[115][143],
reservoir_weight[115][144],
reservoir_weight[115][145],
reservoir_weight[115][146],
reservoir_weight[115][147],
reservoir_weight[115][148],
reservoir_weight[115][149],
reservoir_weight[115][150],
reservoir_weight[115][151],
reservoir_weight[115][152],
reservoir_weight[115][153],
reservoir_weight[115][154],
reservoir_weight[115][155],
reservoir_weight[115][156],
reservoir_weight[115][157],
reservoir_weight[115][158],
reservoir_weight[115][159],
reservoir_weight[115][160],
reservoir_weight[115][161],
reservoir_weight[115][162],
reservoir_weight[115][163],
reservoir_weight[115][164],
reservoir_weight[115][165],
reservoir_weight[115][166],
reservoir_weight[115][167],
reservoir_weight[115][168],
reservoir_weight[115][169],
reservoir_weight[115][170],
reservoir_weight[115][171],
reservoir_weight[115][172],
reservoir_weight[115][173],
reservoir_weight[115][174],
reservoir_weight[115][175],
reservoir_weight[115][176],
reservoir_weight[115][177],
reservoir_weight[115][178],
reservoir_weight[115][179],
reservoir_weight[115][180],
reservoir_weight[115][181],
reservoir_weight[115][182],
reservoir_weight[115][183],
reservoir_weight[115][184],
reservoir_weight[115][185],
reservoir_weight[115][186],
reservoir_weight[115][187],
reservoir_weight[115][188],
reservoir_weight[115][189],
reservoir_weight[115][190],
reservoir_weight[115][191],
reservoir_weight[115][192],
reservoir_weight[115][193],
reservoir_weight[115][194],
reservoir_weight[115][195],
reservoir_weight[115][196],
reservoir_weight[115][197],
reservoir_weight[115][198],
reservoir_weight[115][199]
},
{reservoir_weight[116][0],
reservoir_weight[116][1],
reservoir_weight[116][2],
reservoir_weight[116][3],
reservoir_weight[116][4],
reservoir_weight[116][5],
reservoir_weight[116][6],
reservoir_weight[116][7],
reservoir_weight[116][8],
reservoir_weight[116][9],
reservoir_weight[116][10],
reservoir_weight[116][11],
reservoir_weight[116][12],
reservoir_weight[116][13],
reservoir_weight[116][14],
reservoir_weight[116][15],
reservoir_weight[116][16],
reservoir_weight[116][17],
reservoir_weight[116][18],
reservoir_weight[116][19],
reservoir_weight[116][20],
reservoir_weight[116][21],
reservoir_weight[116][22],
reservoir_weight[116][23],
reservoir_weight[116][24],
reservoir_weight[116][25],
reservoir_weight[116][26],
reservoir_weight[116][27],
reservoir_weight[116][28],
reservoir_weight[116][29],
reservoir_weight[116][30],
reservoir_weight[116][31],
reservoir_weight[116][32],
reservoir_weight[116][33],
reservoir_weight[116][34],
reservoir_weight[116][35],
reservoir_weight[116][36],
reservoir_weight[116][37],
reservoir_weight[116][38],
reservoir_weight[116][39],
reservoir_weight[116][40],
reservoir_weight[116][41],
reservoir_weight[116][42],
reservoir_weight[116][43],
reservoir_weight[116][44],
reservoir_weight[116][45],
reservoir_weight[116][46],
reservoir_weight[116][47],
reservoir_weight[116][48],
reservoir_weight[116][49],
reservoir_weight[116][50],
reservoir_weight[116][51],
reservoir_weight[116][52],
reservoir_weight[116][53],
reservoir_weight[116][54],
reservoir_weight[116][55],
reservoir_weight[116][56],
reservoir_weight[116][57],
reservoir_weight[116][58],
reservoir_weight[116][59],
reservoir_weight[116][60],
reservoir_weight[116][61],
reservoir_weight[116][62],
reservoir_weight[116][63],
reservoir_weight[116][64],
reservoir_weight[116][65],
reservoir_weight[116][66],
reservoir_weight[116][67],
reservoir_weight[116][68],
reservoir_weight[116][69],
reservoir_weight[116][70],
reservoir_weight[116][71],
reservoir_weight[116][72],
reservoir_weight[116][73],
reservoir_weight[116][74],
reservoir_weight[116][75],
reservoir_weight[116][76],
reservoir_weight[116][77],
reservoir_weight[116][78],
reservoir_weight[116][79],
reservoir_weight[116][80],
reservoir_weight[116][81],
reservoir_weight[116][82],
reservoir_weight[116][83],
reservoir_weight[116][84],
reservoir_weight[116][85],
reservoir_weight[116][86],
reservoir_weight[116][87],
reservoir_weight[116][88],
reservoir_weight[116][89],
reservoir_weight[116][90],
reservoir_weight[116][91],
reservoir_weight[116][92],
reservoir_weight[116][93],
reservoir_weight[116][94],
reservoir_weight[116][95],
reservoir_weight[116][96],
reservoir_weight[116][97],
reservoir_weight[116][98],
reservoir_weight[116][99],
reservoir_weight[116][100],
reservoir_weight[116][101],
reservoir_weight[116][102],
reservoir_weight[116][103],
reservoir_weight[116][104],
reservoir_weight[116][105],
reservoir_weight[116][106],
reservoir_weight[116][107],
reservoir_weight[116][108],
reservoir_weight[116][109],
reservoir_weight[116][110],
reservoir_weight[116][111],
reservoir_weight[116][112],
reservoir_weight[116][113],
reservoir_weight[116][114],
reservoir_weight[116][115],
reservoir_weight[116][116],
reservoir_weight[116][117],
reservoir_weight[116][118],
reservoir_weight[116][119],
reservoir_weight[116][120],
reservoir_weight[116][121],
reservoir_weight[116][122],
reservoir_weight[116][123],
reservoir_weight[116][124],
reservoir_weight[116][125],
reservoir_weight[116][126],
reservoir_weight[116][127],
reservoir_weight[116][128],
reservoir_weight[116][129],
reservoir_weight[116][130],
reservoir_weight[116][131],
reservoir_weight[116][132],
reservoir_weight[116][133],
reservoir_weight[116][134],
reservoir_weight[116][135],
reservoir_weight[116][136],
reservoir_weight[116][137],
reservoir_weight[116][138],
reservoir_weight[116][139],
reservoir_weight[116][140],
reservoir_weight[116][141],
reservoir_weight[116][142],
reservoir_weight[116][143],
reservoir_weight[116][144],
reservoir_weight[116][145],
reservoir_weight[116][146],
reservoir_weight[116][147],
reservoir_weight[116][148],
reservoir_weight[116][149],
reservoir_weight[116][150],
reservoir_weight[116][151],
reservoir_weight[116][152],
reservoir_weight[116][153],
reservoir_weight[116][154],
reservoir_weight[116][155],
reservoir_weight[116][156],
reservoir_weight[116][157],
reservoir_weight[116][158],
reservoir_weight[116][159],
reservoir_weight[116][160],
reservoir_weight[116][161],
reservoir_weight[116][162],
reservoir_weight[116][163],
reservoir_weight[116][164],
reservoir_weight[116][165],
reservoir_weight[116][166],
reservoir_weight[116][167],
reservoir_weight[116][168],
reservoir_weight[116][169],
reservoir_weight[116][170],
reservoir_weight[116][171],
reservoir_weight[116][172],
reservoir_weight[116][173],
reservoir_weight[116][174],
reservoir_weight[116][175],
reservoir_weight[116][176],
reservoir_weight[116][177],
reservoir_weight[116][178],
reservoir_weight[116][179],
reservoir_weight[116][180],
reservoir_weight[116][181],
reservoir_weight[116][182],
reservoir_weight[116][183],
reservoir_weight[116][184],
reservoir_weight[116][185],
reservoir_weight[116][186],
reservoir_weight[116][187],
reservoir_weight[116][188],
reservoir_weight[116][189],
reservoir_weight[116][190],
reservoir_weight[116][191],
reservoir_weight[116][192],
reservoir_weight[116][193],
reservoir_weight[116][194],
reservoir_weight[116][195],
reservoir_weight[116][196],
reservoir_weight[116][197],
reservoir_weight[116][198],
reservoir_weight[116][199]
},
{reservoir_weight[117][0],
reservoir_weight[117][1],
reservoir_weight[117][2],
reservoir_weight[117][3],
reservoir_weight[117][4],
reservoir_weight[117][5],
reservoir_weight[117][6],
reservoir_weight[117][7],
reservoir_weight[117][8],
reservoir_weight[117][9],
reservoir_weight[117][10],
reservoir_weight[117][11],
reservoir_weight[117][12],
reservoir_weight[117][13],
reservoir_weight[117][14],
reservoir_weight[117][15],
reservoir_weight[117][16],
reservoir_weight[117][17],
reservoir_weight[117][18],
reservoir_weight[117][19],
reservoir_weight[117][20],
reservoir_weight[117][21],
reservoir_weight[117][22],
reservoir_weight[117][23],
reservoir_weight[117][24],
reservoir_weight[117][25],
reservoir_weight[117][26],
reservoir_weight[117][27],
reservoir_weight[117][28],
reservoir_weight[117][29],
reservoir_weight[117][30],
reservoir_weight[117][31],
reservoir_weight[117][32],
reservoir_weight[117][33],
reservoir_weight[117][34],
reservoir_weight[117][35],
reservoir_weight[117][36],
reservoir_weight[117][37],
reservoir_weight[117][38],
reservoir_weight[117][39],
reservoir_weight[117][40],
reservoir_weight[117][41],
reservoir_weight[117][42],
reservoir_weight[117][43],
reservoir_weight[117][44],
reservoir_weight[117][45],
reservoir_weight[117][46],
reservoir_weight[117][47],
reservoir_weight[117][48],
reservoir_weight[117][49],
reservoir_weight[117][50],
reservoir_weight[117][51],
reservoir_weight[117][52],
reservoir_weight[117][53],
reservoir_weight[117][54],
reservoir_weight[117][55],
reservoir_weight[117][56],
reservoir_weight[117][57],
reservoir_weight[117][58],
reservoir_weight[117][59],
reservoir_weight[117][60],
reservoir_weight[117][61],
reservoir_weight[117][62],
reservoir_weight[117][63],
reservoir_weight[117][64],
reservoir_weight[117][65],
reservoir_weight[117][66],
reservoir_weight[117][67],
reservoir_weight[117][68],
reservoir_weight[117][69],
reservoir_weight[117][70],
reservoir_weight[117][71],
reservoir_weight[117][72],
reservoir_weight[117][73],
reservoir_weight[117][74],
reservoir_weight[117][75],
reservoir_weight[117][76],
reservoir_weight[117][77],
reservoir_weight[117][78],
reservoir_weight[117][79],
reservoir_weight[117][80],
reservoir_weight[117][81],
reservoir_weight[117][82],
reservoir_weight[117][83],
reservoir_weight[117][84],
reservoir_weight[117][85],
reservoir_weight[117][86],
reservoir_weight[117][87],
reservoir_weight[117][88],
reservoir_weight[117][89],
reservoir_weight[117][90],
reservoir_weight[117][91],
reservoir_weight[117][92],
reservoir_weight[117][93],
reservoir_weight[117][94],
reservoir_weight[117][95],
reservoir_weight[117][96],
reservoir_weight[117][97],
reservoir_weight[117][98],
reservoir_weight[117][99],
reservoir_weight[117][100],
reservoir_weight[117][101],
reservoir_weight[117][102],
reservoir_weight[117][103],
reservoir_weight[117][104],
reservoir_weight[117][105],
reservoir_weight[117][106],
reservoir_weight[117][107],
reservoir_weight[117][108],
reservoir_weight[117][109],
reservoir_weight[117][110],
reservoir_weight[117][111],
reservoir_weight[117][112],
reservoir_weight[117][113],
reservoir_weight[117][114],
reservoir_weight[117][115],
reservoir_weight[117][116],
reservoir_weight[117][117],
reservoir_weight[117][118],
reservoir_weight[117][119],
reservoir_weight[117][120],
reservoir_weight[117][121],
reservoir_weight[117][122],
reservoir_weight[117][123],
reservoir_weight[117][124],
reservoir_weight[117][125],
reservoir_weight[117][126],
reservoir_weight[117][127],
reservoir_weight[117][128],
reservoir_weight[117][129],
reservoir_weight[117][130],
reservoir_weight[117][131],
reservoir_weight[117][132],
reservoir_weight[117][133],
reservoir_weight[117][134],
reservoir_weight[117][135],
reservoir_weight[117][136],
reservoir_weight[117][137],
reservoir_weight[117][138],
reservoir_weight[117][139],
reservoir_weight[117][140],
reservoir_weight[117][141],
reservoir_weight[117][142],
reservoir_weight[117][143],
reservoir_weight[117][144],
reservoir_weight[117][145],
reservoir_weight[117][146],
reservoir_weight[117][147],
reservoir_weight[117][148],
reservoir_weight[117][149],
reservoir_weight[117][150],
reservoir_weight[117][151],
reservoir_weight[117][152],
reservoir_weight[117][153],
reservoir_weight[117][154],
reservoir_weight[117][155],
reservoir_weight[117][156],
reservoir_weight[117][157],
reservoir_weight[117][158],
reservoir_weight[117][159],
reservoir_weight[117][160],
reservoir_weight[117][161],
reservoir_weight[117][162],
reservoir_weight[117][163],
reservoir_weight[117][164],
reservoir_weight[117][165],
reservoir_weight[117][166],
reservoir_weight[117][167],
reservoir_weight[117][168],
reservoir_weight[117][169],
reservoir_weight[117][170],
reservoir_weight[117][171],
reservoir_weight[117][172],
reservoir_weight[117][173],
reservoir_weight[117][174],
reservoir_weight[117][175],
reservoir_weight[117][176],
reservoir_weight[117][177],
reservoir_weight[117][178],
reservoir_weight[117][179],
reservoir_weight[117][180],
reservoir_weight[117][181],
reservoir_weight[117][182],
reservoir_weight[117][183],
reservoir_weight[117][184],
reservoir_weight[117][185],
reservoir_weight[117][186],
reservoir_weight[117][187],
reservoir_weight[117][188],
reservoir_weight[117][189],
reservoir_weight[117][190],
reservoir_weight[117][191],
reservoir_weight[117][192],
reservoir_weight[117][193],
reservoir_weight[117][194],
reservoir_weight[117][195],
reservoir_weight[117][196],
reservoir_weight[117][197],
reservoir_weight[117][198],
reservoir_weight[117][199]
},
{reservoir_weight[118][0],
reservoir_weight[118][1],
reservoir_weight[118][2],
reservoir_weight[118][3],
reservoir_weight[118][4],
reservoir_weight[118][5],
reservoir_weight[118][6],
reservoir_weight[118][7],
reservoir_weight[118][8],
reservoir_weight[118][9],
reservoir_weight[118][10],
reservoir_weight[118][11],
reservoir_weight[118][12],
reservoir_weight[118][13],
reservoir_weight[118][14],
reservoir_weight[118][15],
reservoir_weight[118][16],
reservoir_weight[118][17],
reservoir_weight[118][18],
reservoir_weight[118][19],
reservoir_weight[118][20],
reservoir_weight[118][21],
reservoir_weight[118][22],
reservoir_weight[118][23],
reservoir_weight[118][24],
reservoir_weight[118][25],
reservoir_weight[118][26],
reservoir_weight[118][27],
reservoir_weight[118][28],
reservoir_weight[118][29],
reservoir_weight[118][30],
reservoir_weight[118][31],
reservoir_weight[118][32],
reservoir_weight[118][33],
reservoir_weight[118][34],
reservoir_weight[118][35],
reservoir_weight[118][36],
reservoir_weight[118][37],
reservoir_weight[118][38],
reservoir_weight[118][39],
reservoir_weight[118][40],
reservoir_weight[118][41],
reservoir_weight[118][42],
reservoir_weight[118][43],
reservoir_weight[118][44],
reservoir_weight[118][45],
reservoir_weight[118][46],
reservoir_weight[118][47],
reservoir_weight[118][48],
reservoir_weight[118][49],
reservoir_weight[118][50],
reservoir_weight[118][51],
reservoir_weight[118][52],
reservoir_weight[118][53],
reservoir_weight[118][54],
reservoir_weight[118][55],
reservoir_weight[118][56],
reservoir_weight[118][57],
reservoir_weight[118][58],
reservoir_weight[118][59],
reservoir_weight[118][60],
reservoir_weight[118][61],
reservoir_weight[118][62],
reservoir_weight[118][63],
reservoir_weight[118][64],
reservoir_weight[118][65],
reservoir_weight[118][66],
reservoir_weight[118][67],
reservoir_weight[118][68],
reservoir_weight[118][69],
reservoir_weight[118][70],
reservoir_weight[118][71],
reservoir_weight[118][72],
reservoir_weight[118][73],
reservoir_weight[118][74],
reservoir_weight[118][75],
reservoir_weight[118][76],
reservoir_weight[118][77],
reservoir_weight[118][78],
reservoir_weight[118][79],
reservoir_weight[118][80],
reservoir_weight[118][81],
reservoir_weight[118][82],
reservoir_weight[118][83],
reservoir_weight[118][84],
reservoir_weight[118][85],
reservoir_weight[118][86],
reservoir_weight[118][87],
reservoir_weight[118][88],
reservoir_weight[118][89],
reservoir_weight[118][90],
reservoir_weight[118][91],
reservoir_weight[118][92],
reservoir_weight[118][93],
reservoir_weight[118][94],
reservoir_weight[118][95],
reservoir_weight[118][96],
reservoir_weight[118][97],
reservoir_weight[118][98],
reservoir_weight[118][99],
reservoir_weight[118][100],
reservoir_weight[118][101],
reservoir_weight[118][102],
reservoir_weight[118][103],
reservoir_weight[118][104],
reservoir_weight[118][105],
reservoir_weight[118][106],
reservoir_weight[118][107],
reservoir_weight[118][108],
reservoir_weight[118][109],
reservoir_weight[118][110],
reservoir_weight[118][111],
reservoir_weight[118][112],
reservoir_weight[118][113],
reservoir_weight[118][114],
reservoir_weight[118][115],
reservoir_weight[118][116],
reservoir_weight[118][117],
reservoir_weight[118][118],
reservoir_weight[118][119],
reservoir_weight[118][120],
reservoir_weight[118][121],
reservoir_weight[118][122],
reservoir_weight[118][123],
reservoir_weight[118][124],
reservoir_weight[118][125],
reservoir_weight[118][126],
reservoir_weight[118][127],
reservoir_weight[118][128],
reservoir_weight[118][129],
reservoir_weight[118][130],
reservoir_weight[118][131],
reservoir_weight[118][132],
reservoir_weight[118][133],
reservoir_weight[118][134],
reservoir_weight[118][135],
reservoir_weight[118][136],
reservoir_weight[118][137],
reservoir_weight[118][138],
reservoir_weight[118][139],
reservoir_weight[118][140],
reservoir_weight[118][141],
reservoir_weight[118][142],
reservoir_weight[118][143],
reservoir_weight[118][144],
reservoir_weight[118][145],
reservoir_weight[118][146],
reservoir_weight[118][147],
reservoir_weight[118][148],
reservoir_weight[118][149],
reservoir_weight[118][150],
reservoir_weight[118][151],
reservoir_weight[118][152],
reservoir_weight[118][153],
reservoir_weight[118][154],
reservoir_weight[118][155],
reservoir_weight[118][156],
reservoir_weight[118][157],
reservoir_weight[118][158],
reservoir_weight[118][159],
reservoir_weight[118][160],
reservoir_weight[118][161],
reservoir_weight[118][162],
reservoir_weight[118][163],
reservoir_weight[118][164],
reservoir_weight[118][165],
reservoir_weight[118][166],
reservoir_weight[118][167],
reservoir_weight[118][168],
reservoir_weight[118][169],
reservoir_weight[118][170],
reservoir_weight[118][171],
reservoir_weight[118][172],
reservoir_weight[118][173],
reservoir_weight[118][174],
reservoir_weight[118][175],
reservoir_weight[118][176],
reservoir_weight[118][177],
reservoir_weight[118][178],
reservoir_weight[118][179],
reservoir_weight[118][180],
reservoir_weight[118][181],
reservoir_weight[118][182],
reservoir_weight[118][183],
reservoir_weight[118][184],
reservoir_weight[118][185],
reservoir_weight[118][186],
reservoir_weight[118][187],
reservoir_weight[118][188],
reservoir_weight[118][189],
reservoir_weight[118][190],
reservoir_weight[118][191],
reservoir_weight[118][192],
reservoir_weight[118][193],
reservoir_weight[118][194],
reservoir_weight[118][195],
reservoir_weight[118][196],
reservoir_weight[118][197],
reservoir_weight[118][198],
reservoir_weight[118][199]
},
{reservoir_weight[119][0],
reservoir_weight[119][1],
reservoir_weight[119][2],
reservoir_weight[119][3],
reservoir_weight[119][4],
reservoir_weight[119][5],
reservoir_weight[119][6],
reservoir_weight[119][7],
reservoir_weight[119][8],
reservoir_weight[119][9],
reservoir_weight[119][10],
reservoir_weight[119][11],
reservoir_weight[119][12],
reservoir_weight[119][13],
reservoir_weight[119][14],
reservoir_weight[119][15],
reservoir_weight[119][16],
reservoir_weight[119][17],
reservoir_weight[119][18],
reservoir_weight[119][19],
reservoir_weight[119][20],
reservoir_weight[119][21],
reservoir_weight[119][22],
reservoir_weight[119][23],
reservoir_weight[119][24],
reservoir_weight[119][25],
reservoir_weight[119][26],
reservoir_weight[119][27],
reservoir_weight[119][28],
reservoir_weight[119][29],
reservoir_weight[119][30],
reservoir_weight[119][31],
reservoir_weight[119][32],
reservoir_weight[119][33],
reservoir_weight[119][34],
reservoir_weight[119][35],
reservoir_weight[119][36],
reservoir_weight[119][37],
reservoir_weight[119][38],
reservoir_weight[119][39],
reservoir_weight[119][40],
reservoir_weight[119][41],
reservoir_weight[119][42],
reservoir_weight[119][43],
reservoir_weight[119][44],
reservoir_weight[119][45],
reservoir_weight[119][46],
reservoir_weight[119][47],
reservoir_weight[119][48],
reservoir_weight[119][49],
reservoir_weight[119][50],
reservoir_weight[119][51],
reservoir_weight[119][52],
reservoir_weight[119][53],
reservoir_weight[119][54],
reservoir_weight[119][55],
reservoir_weight[119][56],
reservoir_weight[119][57],
reservoir_weight[119][58],
reservoir_weight[119][59],
reservoir_weight[119][60],
reservoir_weight[119][61],
reservoir_weight[119][62],
reservoir_weight[119][63],
reservoir_weight[119][64],
reservoir_weight[119][65],
reservoir_weight[119][66],
reservoir_weight[119][67],
reservoir_weight[119][68],
reservoir_weight[119][69],
reservoir_weight[119][70],
reservoir_weight[119][71],
reservoir_weight[119][72],
reservoir_weight[119][73],
reservoir_weight[119][74],
reservoir_weight[119][75],
reservoir_weight[119][76],
reservoir_weight[119][77],
reservoir_weight[119][78],
reservoir_weight[119][79],
reservoir_weight[119][80],
reservoir_weight[119][81],
reservoir_weight[119][82],
reservoir_weight[119][83],
reservoir_weight[119][84],
reservoir_weight[119][85],
reservoir_weight[119][86],
reservoir_weight[119][87],
reservoir_weight[119][88],
reservoir_weight[119][89],
reservoir_weight[119][90],
reservoir_weight[119][91],
reservoir_weight[119][92],
reservoir_weight[119][93],
reservoir_weight[119][94],
reservoir_weight[119][95],
reservoir_weight[119][96],
reservoir_weight[119][97],
reservoir_weight[119][98],
reservoir_weight[119][99],
reservoir_weight[119][100],
reservoir_weight[119][101],
reservoir_weight[119][102],
reservoir_weight[119][103],
reservoir_weight[119][104],
reservoir_weight[119][105],
reservoir_weight[119][106],
reservoir_weight[119][107],
reservoir_weight[119][108],
reservoir_weight[119][109],
reservoir_weight[119][110],
reservoir_weight[119][111],
reservoir_weight[119][112],
reservoir_weight[119][113],
reservoir_weight[119][114],
reservoir_weight[119][115],
reservoir_weight[119][116],
reservoir_weight[119][117],
reservoir_weight[119][118],
reservoir_weight[119][119],
reservoir_weight[119][120],
reservoir_weight[119][121],
reservoir_weight[119][122],
reservoir_weight[119][123],
reservoir_weight[119][124],
reservoir_weight[119][125],
reservoir_weight[119][126],
reservoir_weight[119][127],
reservoir_weight[119][128],
reservoir_weight[119][129],
reservoir_weight[119][130],
reservoir_weight[119][131],
reservoir_weight[119][132],
reservoir_weight[119][133],
reservoir_weight[119][134],
reservoir_weight[119][135],
reservoir_weight[119][136],
reservoir_weight[119][137],
reservoir_weight[119][138],
reservoir_weight[119][139],
reservoir_weight[119][140],
reservoir_weight[119][141],
reservoir_weight[119][142],
reservoir_weight[119][143],
reservoir_weight[119][144],
reservoir_weight[119][145],
reservoir_weight[119][146],
reservoir_weight[119][147],
reservoir_weight[119][148],
reservoir_weight[119][149],
reservoir_weight[119][150],
reservoir_weight[119][151],
reservoir_weight[119][152],
reservoir_weight[119][153],
reservoir_weight[119][154],
reservoir_weight[119][155],
reservoir_weight[119][156],
reservoir_weight[119][157],
reservoir_weight[119][158],
reservoir_weight[119][159],
reservoir_weight[119][160],
reservoir_weight[119][161],
reservoir_weight[119][162],
reservoir_weight[119][163],
reservoir_weight[119][164],
reservoir_weight[119][165],
reservoir_weight[119][166],
reservoir_weight[119][167],
reservoir_weight[119][168],
reservoir_weight[119][169],
reservoir_weight[119][170],
reservoir_weight[119][171],
reservoir_weight[119][172],
reservoir_weight[119][173],
reservoir_weight[119][174],
reservoir_weight[119][175],
reservoir_weight[119][176],
reservoir_weight[119][177],
reservoir_weight[119][178],
reservoir_weight[119][179],
reservoir_weight[119][180],
reservoir_weight[119][181],
reservoir_weight[119][182],
reservoir_weight[119][183],
reservoir_weight[119][184],
reservoir_weight[119][185],
reservoir_weight[119][186],
reservoir_weight[119][187],
reservoir_weight[119][188],
reservoir_weight[119][189],
reservoir_weight[119][190],
reservoir_weight[119][191],
reservoir_weight[119][192],
reservoir_weight[119][193],
reservoir_weight[119][194],
reservoir_weight[119][195],
reservoir_weight[119][196],
reservoir_weight[119][197],
reservoir_weight[119][198],
reservoir_weight[119][199]
},
{reservoir_weight[120][0],
reservoir_weight[120][1],
reservoir_weight[120][2],
reservoir_weight[120][3],
reservoir_weight[120][4],
reservoir_weight[120][5],
reservoir_weight[120][6],
reservoir_weight[120][7],
reservoir_weight[120][8],
reservoir_weight[120][9],
reservoir_weight[120][10],
reservoir_weight[120][11],
reservoir_weight[120][12],
reservoir_weight[120][13],
reservoir_weight[120][14],
reservoir_weight[120][15],
reservoir_weight[120][16],
reservoir_weight[120][17],
reservoir_weight[120][18],
reservoir_weight[120][19],
reservoir_weight[120][20],
reservoir_weight[120][21],
reservoir_weight[120][22],
reservoir_weight[120][23],
reservoir_weight[120][24],
reservoir_weight[120][25],
reservoir_weight[120][26],
reservoir_weight[120][27],
reservoir_weight[120][28],
reservoir_weight[120][29],
reservoir_weight[120][30],
reservoir_weight[120][31],
reservoir_weight[120][32],
reservoir_weight[120][33],
reservoir_weight[120][34],
reservoir_weight[120][35],
reservoir_weight[120][36],
reservoir_weight[120][37],
reservoir_weight[120][38],
reservoir_weight[120][39],
reservoir_weight[120][40],
reservoir_weight[120][41],
reservoir_weight[120][42],
reservoir_weight[120][43],
reservoir_weight[120][44],
reservoir_weight[120][45],
reservoir_weight[120][46],
reservoir_weight[120][47],
reservoir_weight[120][48],
reservoir_weight[120][49],
reservoir_weight[120][50],
reservoir_weight[120][51],
reservoir_weight[120][52],
reservoir_weight[120][53],
reservoir_weight[120][54],
reservoir_weight[120][55],
reservoir_weight[120][56],
reservoir_weight[120][57],
reservoir_weight[120][58],
reservoir_weight[120][59],
reservoir_weight[120][60],
reservoir_weight[120][61],
reservoir_weight[120][62],
reservoir_weight[120][63],
reservoir_weight[120][64],
reservoir_weight[120][65],
reservoir_weight[120][66],
reservoir_weight[120][67],
reservoir_weight[120][68],
reservoir_weight[120][69],
reservoir_weight[120][70],
reservoir_weight[120][71],
reservoir_weight[120][72],
reservoir_weight[120][73],
reservoir_weight[120][74],
reservoir_weight[120][75],
reservoir_weight[120][76],
reservoir_weight[120][77],
reservoir_weight[120][78],
reservoir_weight[120][79],
reservoir_weight[120][80],
reservoir_weight[120][81],
reservoir_weight[120][82],
reservoir_weight[120][83],
reservoir_weight[120][84],
reservoir_weight[120][85],
reservoir_weight[120][86],
reservoir_weight[120][87],
reservoir_weight[120][88],
reservoir_weight[120][89],
reservoir_weight[120][90],
reservoir_weight[120][91],
reservoir_weight[120][92],
reservoir_weight[120][93],
reservoir_weight[120][94],
reservoir_weight[120][95],
reservoir_weight[120][96],
reservoir_weight[120][97],
reservoir_weight[120][98],
reservoir_weight[120][99],
reservoir_weight[120][100],
reservoir_weight[120][101],
reservoir_weight[120][102],
reservoir_weight[120][103],
reservoir_weight[120][104],
reservoir_weight[120][105],
reservoir_weight[120][106],
reservoir_weight[120][107],
reservoir_weight[120][108],
reservoir_weight[120][109],
reservoir_weight[120][110],
reservoir_weight[120][111],
reservoir_weight[120][112],
reservoir_weight[120][113],
reservoir_weight[120][114],
reservoir_weight[120][115],
reservoir_weight[120][116],
reservoir_weight[120][117],
reservoir_weight[120][118],
reservoir_weight[120][119],
reservoir_weight[120][120],
reservoir_weight[120][121],
reservoir_weight[120][122],
reservoir_weight[120][123],
reservoir_weight[120][124],
reservoir_weight[120][125],
reservoir_weight[120][126],
reservoir_weight[120][127],
reservoir_weight[120][128],
reservoir_weight[120][129],
reservoir_weight[120][130],
reservoir_weight[120][131],
reservoir_weight[120][132],
reservoir_weight[120][133],
reservoir_weight[120][134],
reservoir_weight[120][135],
reservoir_weight[120][136],
reservoir_weight[120][137],
reservoir_weight[120][138],
reservoir_weight[120][139],
reservoir_weight[120][140],
reservoir_weight[120][141],
reservoir_weight[120][142],
reservoir_weight[120][143],
reservoir_weight[120][144],
reservoir_weight[120][145],
reservoir_weight[120][146],
reservoir_weight[120][147],
reservoir_weight[120][148],
reservoir_weight[120][149],
reservoir_weight[120][150],
reservoir_weight[120][151],
reservoir_weight[120][152],
reservoir_weight[120][153],
reservoir_weight[120][154],
reservoir_weight[120][155],
reservoir_weight[120][156],
reservoir_weight[120][157],
reservoir_weight[120][158],
reservoir_weight[120][159],
reservoir_weight[120][160],
reservoir_weight[120][161],
reservoir_weight[120][162],
reservoir_weight[120][163],
reservoir_weight[120][164],
reservoir_weight[120][165],
reservoir_weight[120][166],
reservoir_weight[120][167],
reservoir_weight[120][168],
reservoir_weight[120][169],
reservoir_weight[120][170],
reservoir_weight[120][171],
reservoir_weight[120][172],
reservoir_weight[120][173],
reservoir_weight[120][174],
reservoir_weight[120][175],
reservoir_weight[120][176],
reservoir_weight[120][177],
reservoir_weight[120][178],
reservoir_weight[120][179],
reservoir_weight[120][180],
reservoir_weight[120][181],
reservoir_weight[120][182],
reservoir_weight[120][183],
reservoir_weight[120][184],
reservoir_weight[120][185],
reservoir_weight[120][186],
reservoir_weight[120][187],
reservoir_weight[120][188],
reservoir_weight[120][189],
reservoir_weight[120][190],
reservoir_weight[120][191],
reservoir_weight[120][192],
reservoir_weight[120][193],
reservoir_weight[120][194],
reservoir_weight[120][195],
reservoir_weight[120][196],
reservoir_weight[120][197],
reservoir_weight[120][198],
reservoir_weight[120][199]
},
{reservoir_weight[121][0],
reservoir_weight[121][1],
reservoir_weight[121][2],
reservoir_weight[121][3],
reservoir_weight[121][4],
reservoir_weight[121][5],
reservoir_weight[121][6],
reservoir_weight[121][7],
reservoir_weight[121][8],
reservoir_weight[121][9],
reservoir_weight[121][10],
reservoir_weight[121][11],
reservoir_weight[121][12],
reservoir_weight[121][13],
reservoir_weight[121][14],
reservoir_weight[121][15],
reservoir_weight[121][16],
reservoir_weight[121][17],
reservoir_weight[121][18],
reservoir_weight[121][19],
reservoir_weight[121][20],
reservoir_weight[121][21],
reservoir_weight[121][22],
reservoir_weight[121][23],
reservoir_weight[121][24],
reservoir_weight[121][25],
reservoir_weight[121][26],
reservoir_weight[121][27],
reservoir_weight[121][28],
reservoir_weight[121][29],
reservoir_weight[121][30],
reservoir_weight[121][31],
reservoir_weight[121][32],
reservoir_weight[121][33],
reservoir_weight[121][34],
reservoir_weight[121][35],
reservoir_weight[121][36],
reservoir_weight[121][37],
reservoir_weight[121][38],
reservoir_weight[121][39],
reservoir_weight[121][40],
reservoir_weight[121][41],
reservoir_weight[121][42],
reservoir_weight[121][43],
reservoir_weight[121][44],
reservoir_weight[121][45],
reservoir_weight[121][46],
reservoir_weight[121][47],
reservoir_weight[121][48],
reservoir_weight[121][49],
reservoir_weight[121][50],
reservoir_weight[121][51],
reservoir_weight[121][52],
reservoir_weight[121][53],
reservoir_weight[121][54],
reservoir_weight[121][55],
reservoir_weight[121][56],
reservoir_weight[121][57],
reservoir_weight[121][58],
reservoir_weight[121][59],
reservoir_weight[121][60],
reservoir_weight[121][61],
reservoir_weight[121][62],
reservoir_weight[121][63],
reservoir_weight[121][64],
reservoir_weight[121][65],
reservoir_weight[121][66],
reservoir_weight[121][67],
reservoir_weight[121][68],
reservoir_weight[121][69],
reservoir_weight[121][70],
reservoir_weight[121][71],
reservoir_weight[121][72],
reservoir_weight[121][73],
reservoir_weight[121][74],
reservoir_weight[121][75],
reservoir_weight[121][76],
reservoir_weight[121][77],
reservoir_weight[121][78],
reservoir_weight[121][79],
reservoir_weight[121][80],
reservoir_weight[121][81],
reservoir_weight[121][82],
reservoir_weight[121][83],
reservoir_weight[121][84],
reservoir_weight[121][85],
reservoir_weight[121][86],
reservoir_weight[121][87],
reservoir_weight[121][88],
reservoir_weight[121][89],
reservoir_weight[121][90],
reservoir_weight[121][91],
reservoir_weight[121][92],
reservoir_weight[121][93],
reservoir_weight[121][94],
reservoir_weight[121][95],
reservoir_weight[121][96],
reservoir_weight[121][97],
reservoir_weight[121][98],
reservoir_weight[121][99],
reservoir_weight[121][100],
reservoir_weight[121][101],
reservoir_weight[121][102],
reservoir_weight[121][103],
reservoir_weight[121][104],
reservoir_weight[121][105],
reservoir_weight[121][106],
reservoir_weight[121][107],
reservoir_weight[121][108],
reservoir_weight[121][109],
reservoir_weight[121][110],
reservoir_weight[121][111],
reservoir_weight[121][112],
reservoir_weight[121][113],
reservoir_weight[121][114],
reservoir_weight[121][115],
reservoir_weight[121][116],
reservoir_weight[121][117],
reservoir_weight[121][118],
reservoir_weight[121][119],
reservoir_weight[121][120],
reservoir_weight[121][121],
reservoir_weight[121][122],
reservoir_weight[121][123],
reservoir_weight[121][124],
reservoir_weight[121][125],
reservoir_weight[121][126],
reservoir_weight[121][127],
reservoir_weight[121][128],
reservoir_weight[121][129],
reservoir_weight[121][130],
reservoir_weight[121][131],
reservoir_weight[121][132],
reservoir_weight[121][133],
reservoir_weight[121][134],
reservoir_weight[121][135],
reservoir_weight[121][136],
reservoir_weight[121][137],
reservoir_weight[121][138],
reservoir_weight[121][139],
reservoir_weight[121][140],
reservoir_weight[121][141],
reservoir_weight[121][142],
reservoir_weight[121][143],
reservoir_weight[121][144],
reservoir_weight[121][145],
reservoir_weight[121][146],
reservoir_weight[121][147],
reservoir_weight[121][148],
reservoir_weight[121][149],
reservoir_weight[121][150],
reservoir_weight[121][151],
reservoir_weight[121][152],
reservoir_weight[121][153],
reservoir_weight[121][154],
reservoir_weight[121][155],
reservoir_weight[121][156],
reservoir_weight[121][157],
reservoir_weight[121][158],
reservoir_weight[121][159],
reservoir_weight[121][160],
reservoir_weight[121][161],
reservoir_weight[121][162],
reservoir_weight[121][163],
reservoir_weight[121][164],
reservoir_weight[121][165],
reservoir_weight[121][166],
reservoir_weight[121][167],
reservoir_weight[121][168],
reservoir_weight[121][169],
reservoir_weight[121][170],
reservoir_weight[121][171],
reservoir_weight[121][172],
reservoir_weight[121][173],
reservoir_weight[121][174],
reservoir_weight[121][175],
reservoir_weight[121][176],
reservoir_weight[121][177],
reservoir_weight[121][178],
reservoir_weight[121][179],
reservoir_weight[121][180],
reservoir_weight[121][181],
reservoir_weight[121][182],
reservoir_weight[121][183],
reservoir_weight[121][184],
reservoir_weight[121][185],
reservoir_weight[121][186],
reservoir_weight[121][187],
reservoir_weight[121][188],
reservoir_weight[121][189],
reservoir_weight[121][190],
reservoir_weight[121][191],
reservoir_weight[121][192],
reservoir_weight[121][193],
reservoir_weight[121][194],
reservoir_weight[121][195],
reservoir_weight[121][196],
reservoir_weight[121][197],
reservoir_weight[121][198],
reservoir_weight[121][199]
},
{reservoir_weight[122][0],
reservoir_weight[122][1],
reservoir_weight[122][2],
reservoir_weight[122][3],
reservoir_weight[122][4],
reservoir_weight[122][5],
reservoir_weight[122][6],
reservoir_weight[122][7],
reservoir_weight[122][8],
reservoir_weight[122][9],
reservoir_weight[122][10],
reservoir_weight[122][11],
reservoir_weight[122][12],
reservoir_weight[122][13],
reservoir_weight[122][14],
reservoir_weight[122][15],
reservoir_weight[122][16],
reservoir_weight[122][17],
reservoir_weight[122][18],
reservoir_weight[122][19],
reservoir_weight[122][20],
reservoir_weight[122][21],
reservoir_weight[122][22],
reservoir_weight[122][23],
reservoir_weight[122][24],
reservoir_weight[122][25],
reservoir_weight[122][26],
reservoir_weight[122][27],
reservoir_weight[122][28],
reservoir_weight[122][29],
reservoir_weight[122][30],
reservoir_weight[122][31],
reservoir_weight[122][32],
reservoir_weight[122][33],
reservoir_weight[122][34],
reservoir_weight[122][35],
reservoir_weight[122][36],
reservoir_weight[122][37],
reservoir_weight[122][38],
reservoir_weight[122][39],
reservoir_weight[122][40],
reservoir_weight[122][41],
reservoir_weight[122][42],
reservoir_weight[122][43],
reservoir_weight[122][44],
reservoir_weight[122][45],
reservoir_weight[122][46],
reservoir_weight[122][47],
reservoir_weight[122][48],
reservoir_weight[122][49],
reservoir_weight[122][50],
reservoir_weight[122][51],
reservoir_weight[122][52],
reservoir_weight[122][53],
reservoir_weight[122][54],
reservoir_weight[122][55],
reservoir_weight[122][56],
reservoir_weight[122][57],
reservoir_weight[122][58],
reservoir_weight[122][59],
reservoir_weight[122][60],
reservoir_weight[122][61],
reservoir_weight[122][62],
reservoir_weight[122][63],
reservoir_weight[122][64],
reservoir_weight[122][65],
reservoir_weight[122][66],
reservoir_weight[122][67],
reservoir_weight[122][68],
reservoir_weight[122][69],
reservoir_weight[122][70],
reservoir_weight[122][71],
reservoir_weight[122][72],
reservoir_weight[122][73],
reservoir_weight[122][74],
reservoir_weight[122][75],
reservoir_weight[122][76],
reservoir_weight[122][77],
reservoir_weight[122][78],
reservoir_weight[122][79],
reservoir_weight[122][80],
reservoir_weight[122][81],
reservoir_weight[122][82],
reservoir_weight[122][83],
reservoir_weight[122][84],
reservoir_weight[122][85],
reservoir_weight[122][86],
reservoir_weight[122][87],
reservoir_weight[122][88],
reservoir_weight[122][89],
reservoir_weight[122][90],
reservoir_weight[122][91],
reservoir_weight[122][92],
reservoir_weight[122][93],
reservoir_weight[122][94],
reservoir_weight[122][95],
reservoir_weight[122][96],
reservoir_weight[122][97],
reservoir_weight[122][98],
reservoir_weight[122][99],
reservoir_weight[122][100],
reservoir_weight[122][101],
reservoir_weight[122][102],
reservoir_weight[122][103],
reservoir_weight[122][104],
reservoir_weight[122][105],
reservoir_weight[122][106],
reservoir_weight[122][107],
reservoir_weight[122][108],
reservoir_weight[122][109],
reservoir_weight[122][110],
reservoir_weight[122][111],
reservoir_weight[122][112],
reservoir_weight[122][113],
reservoir_weight[122][114],
reservoir_weight[122][115],
reservoir_weight[122][116],
reservoir_weight[122][117],
reservoir_weight[122][118],
reservoir_weight[122][119],
reservoir_weight[122][120],
reservoir_weight[122][121],
reservoir_weight[122][122],
reservoir_weight[122][123],
reservoir_weight[122][124],
reservoir_weight[122][125],
reservoir_weight[122][126],
reservoir_weight[122][127],
reservoir_weight[122][128],
reservoir_weight[122][129],
reservoir_weight[122][130],
reservoir_weight[122][131],
reservoir_weight[122][132],
reservoir_weight[122][133],
reservoir_weight[122][134],
reservoir_weight[122][135],
reservoir_weight[122][136],
reservoir_weight[122][137],
reservoir_weight[122][138],
reservoir_weight[122][139],
reservoir_weight[122][140],
reservoir_weight[122][141],
reservoir_weight[122][142],
reservoir_weight[122][143],
reservoir_weight[122][144],
reservoir_weight[122][145],
reservoir_weight[122][146],
reservoir_weight[122][147],
reservoir_weight[122][148],
reservoir_weight[122][149],
reservoir_weight[122][150],
reservoir_weight[122][151],
reservoir_weight[122][152],
reservoir_weight[122][153],
reservoir_weight[122][154],
reservoir_weight[122][155],
reservoir_weight[122][156],
reservoir_weight[122][157],
reservoir_weight[122][158],
reservoir_weight[122][159],
reservoir_weight[122][160],
reservoir_weight[122][161],
reservoir_weight[122][162],
reservoir_weight[122][163],
reservoir_weight[122][164],
reservoir_weight[122][165],
reservoir_weight[122][166],
reservoir_weight[122][167],
reservoir_weight[122][168],
reservoir_weight[122][169],
reservoir_weight[122][170],
reservoir_weight[122][171],
reservoir_weight[122][172],
reservoir_weight[122][173],
reservoir_weight[122][174],
reservoir_weight[122][175],
reservoir_weight[122][176],
reservoir_weight[122][177],
reservoir_weight[122][178],
reservoir_weight[122][179],
reservoir_weight[122][180],
reservoir_weight[122][181],
reservoir_weight[122][182],
reservoir_weight[122][183],
reservoir_weight[122][184],
reservoir_weight[122][185],
reservoir_weight[122][186],
reservoir_weight[122][187],
reservoir_weight[122][188],
reservoir_weight[122][189],
reservoir_weight[122][190],
reservoir_weight[122][191],
reservoir_weight[122][192],
reservoir_weight[122][193],
reservoir_weight[122][194],
reservoir_weight[122][195],
reservoir_weight[122][196],
reservoir_weight[122][197],
reservoir_weight[122][198],
reservoir_weight[122][199]
},
{reservoir_weight[123][0],
reservoir_weight[123][1],
reservoir_weight[123][2],
reservoir_weight[123][3],
reservoir_weight[123][4],
reservoir_weight[123][5],
reservoir_weight[123][6],
reservoir_weight[123][7],
reservoir_weight[123][8],
reservoir_weight[123][9],
reservoir_weight[123][10],
reservoir_weight[123][11],
reservoir_weight[123][12],
reservoir_weight[123][13],
reservoir_weight[123][14],
reservoir_weight[123][15],
reservoir_weight[123][16],
reservoir_weight[123][17],
reservoir_weight[123][18],
reservoir_weight[123][19],
reservoir_weight[123][20],
reservoir_weight[123][21],
reservoir_weight[123][22],
reservoir_weight[123][23],
reservoir_weight[123][24],
reservoir_weight[123][25],
reservoir_weight[123][26],
reservoir_weight[123][27],
reservoir_weight[123][28],
reservoir_weight[123][29],
reservoir_weight[123][30],
reservoir_weight[123][31],
reservoir_weight[123][32],
reservoir_weight[123][33],
reservoir_weight[123][34],
reservoir_weight[123][35],
reservoir_weight[123][36],
reservoir_weight[123][37],
reservoir_weight[123][38],
reservoir_weight[123][39],
reservoir_weight[123][40],
reservoir_weight[123][41],
reservoir_weight[123][42],
reservoir_weight[123][43],
reservoir_weight[123][44],
reservoir_weight[123][45],
reservoir_weight[123][46],
reservoir_weight[123][47],
reservoir_weight[123][48],
reservoir_weight[123][49],
reservoir_weight[123][50],
reservoir_weight[123][51],
reservoir_weight[123][52],
reservoir_weight[123][53],
reservoir_weight[123][54],
reservoir_weight[123][55],
reservoir_weight[123][56],
reservoir_weight[123][57],
reservoir_weight[123][58],
reservoir_weight[123][59],
reservoir_weight[123][60],
reservoir_weight[123][61],
reservoir_weight[123][62],
reservoir_weight[123][63],
reservoir_weight[123][64],
reservoir_weight[123][65],
reservoir_weight[123][66],
reservoir_weight[123][67],
reservoir_weight[123][68],
reservoir_weight[123][69],
reservoir_weight[123][70],
reservoir_weight[123][71],
reservoir_weight[123][72],
reservoir_weight[123][73],
reservoir_weight[123][74],
reservoir_weight[123][75],
reservoir_weight[123][76],
reservoir_weight[123][77],
reservoir_weight[123][78],
reservoir_weight[123][79],
reservoir_weight[123][80],
reservoir_weight[123][81],
reservoir_weight[123][82],
reservoir_weight[123][83],
reservoir_weight[123][84],
reservoir_weight[123][85],
reservoir_weight[123][86],
reservoir_weight[123][87],
reservoir_weight[123][88],
reservoir_weight[123][89],
reservoir_weight[123][90],
reservoir_weight[123][91],
reservoir_weight[123][92],
reservoir_weight[123][93],
reservoir_weight[123][94],
reservoir_weight[123][95],
reservoir_weight[123][96],
reservoir_weight[123][97],
reservoir_weight[123][98],
reservoir_weight[123][99],
reservoir_weight[123][100],
reservoir_weight[123][101],
reservoir_weight[123][102],
reservoir_weight[123][103],
reservoir_weight[123][104],
reservoir_weight[123][105],
reservoir_weight[123][106],
reservoir_weight[123][107],
reservoir_weight[123][108],
reservoir_weight[123][109],
reservoir_weight[123][110],
reservoir_weight[123][111],
reservoir_weight[123][112],
reservoir_weight[123][113],
reservoir_weight[123][114],
reservoir_weight[123][115],
reservoir_weight[123][116],
reservoir_weight[123][117],
reservoir_weight[123][118],
reservoir_weight[123][119],
reservoir_weight[123][120],
reservoir_weight[123][121],
reservoir_weight[123][122],
reservoir_weight[123][123],
reservoir_weight[123][124],
reservoir_weight[123][125],
reservoir_weight[123][126],
reservoir_weight[123][127],
reservoir_weight[123][128],
reservoir_weight[123][129],
reservoir_weight[123][130],
reservoir_weight[123][131],
reservoir_weight[123][132],
reservoir_weight[123][133],
reservoir_weight[123][134],
reservoir_weight[123][135],
reservoir_weight[123][136],
reservoir_weight[123][137],
reservoir_weight[123][138],
reservoir_weight[123][139],
reservoir_weight[123][140],
reservoir_weight[123][141],
reservoir_weight[123][142],
reservoir_weight[123][143],
reservoir_weight[123][144],
reservoir_weight[123][145],
reservoir_weight[123][146],
reservoir_weight[123][147],
reservoir_weight[123][148],
reservoir_weight[123][149],
reservoir_weight[123][150],
reservoir_weight[123][151],
reservoir_weight[123][152],
reservoir_weight[123][153],
reservoir_weight[123][154],
reservoir_weight[123][155],
reservoir_weight[123][156],
reservoir_weight[123][157],
reservoir_weight[123][158],
reservoir_weight[123][159],
reservoir_weight[123][160],
reservoir_weight[123][161],
reservoir_weight[123][162],
reservoir_weight[123][163],
reservoir_weight[123][164],
reservoir_weight[123][165],
reservoir_weight[123][166],
reservoir_weight[123][167],
reservoir_weight[123][168],
reservoir_weight[123][169],
reservoir_weight[123][170],
reservoir_weight[123][171],
reservoir_weight[123][172],
reservoir_weight[123][173],
reservoir_weight[123][174],
reservoir_weight[123][175],
reservoir_weight[123][176],
reservoir_weight[123][177],
reservoir_weight[123][178],
reservoir_weight[123][179],
reservoir_weight[123][180],
reservoir_weight[123][181],
reservoir_weight[123][182],
reservoir_weight[123][183],
reservoir_weight[123][184],
reservoir_weight[123][185],
reservoir_weight[123][186],
reservoir_weight[123][187],
reservoir_weight[123][188],
reservoir_weight[123][189],
reservoir_weight[123][190],
reservoir_weight[123][191],
reservoir_weight[123][192],
reservoir_weight[123][193],
reservoir_weight[123][194],
reservoir_weight[123][195],
reservoir_weight[123][196],
reservoir_weight[123][197],
reservoir_weight[123][198],
reservoir_weight[123][199]
},
{reservoir_weight[124][0],
reservoir_weight[124][1],
reservoir_weight[124][2],
reservoir_weight[124][3],
reservoir_weight[124][4],
reservoir_weight[124][5],
reservoir_weight[124][6],
reservoir_weight[124][7],
reservoir_weight[124][8],
reservoir_weight[124][9],
reservoir_weight[124][10],
reservoir_weight[124][11],
reservoir_weight[124][12],
reservoir_weight[124][13],
reservoir_weight[124][14],
reservoir_weight[124][15],
reservoir_weight[124][16],
reservoir_weight[124][17],
reservoir_weight[124][18],
reservoir_weight[124][19],
reservoir_weight[124][20],
reservoir_weight[124][21],
reservoir_weight[124][22],
reservoir_weight[124][23],
reservoir_weight[124][24],
reservoir_weight[124][25],
reservoir_weight[124][26],
reservoir_weight[124][27],
reservoir_weight[124][28],
reservoir_weight[124][29],
reservoir_weight[124][30],
reservoir_weight[124][31],
reservoir_weight[124][32],
reservoir_weight[124][33],
reservoir_weight[124][34],
reservoir_weight[124][35],
reservoir_weight[124][36],
reservoir_weight[124][37],
reservoir_weight[124][38],
reservoir_weight[124][39],
reservoir_weight[124][40],
reservoir_weight[124][41],
reservoir_weight[124][42],
reservoir_weight[124][43],
reservoir_weight[124][44],
reservoir_weight[124][45],
reservoir_weight[124][46],
reservoir_weight[124][47],
reservoir_weight[124][48],
reservoir_weight[124][49],
reservoir_weight[124][50],
reservoir_weight[124][51],
reservoir_weight[124][52],
reservoir_weight[124][53],
reservoir_weight[124][54],
reservoir_weight[124][55],
reservoir_weight[124][56],
reservoir_weight[124][57],
reservoir_weight[124][58],
reservoir_weight[124][59],
reservoir_weight[124][60],
reservoir_weight[124][61],
reservoir_weight[124][62],
reservoir_weight[124][63],
reservoir_weight[124][64],
reservoir_weight[124][65],
reservoir_weight[124][66],
reservoir_weight[124][67],
reservoir_weight[124][68],
reservoir_weight[124][69],
reservoir_weight[124][70],
reservoir_weight[124][71],
reservoir_weight[124][72],
reservoir_weight[124][73],
reservoir_weight[124][74],
reservoir_weight[124][75],
reservoir_weight[124][76],
reservoir_weight[124][77],
reservoir_weight[124][78],
reservoir_weight[124][79],
reservoir_weight[124][80],
reservoir_weight[124][81],
reservoir_weight[124][82],
reservoir_weight[124][83],
reservoir_weight[124][84],
reservoir_weight[124][85],
reservoir_weight[124][86],
reservoir_weight[124][87],
reservoir_weight[124][88],
reservoir_weight[124][89],
reservoir_weight[124][90],
reservoir_weight[124][91],
reservoir_weight[124][92],
reservoir_weight[124][93],
reservoir_weight[124][94],
reservoir_weight[124][95],
reservoir_weight[124][96],
reservoir_weight[124][97],
reservoir_weight[124][98],
reservoir_weight[124][99],
reservoir_weight[124][100],
reservoir_weight[124][101],
reservoir_weight[124][102],
reservoir_weight[124][103],
reservoir_weight[124][104],
reservoir_weight[124][105],
reservoir_weight[124][106],
reservoir_weight[124][107],
reservoir_weight[124][108],
reservoir_weight[124][109],
reservoir_weight[124][110],
reservoir_weight[124][111],
reservoir_weight[124][112],
reservoir_weight[124][113],
reservoir_weight[124][114],
reservoir_weight[124][115],
reservoir_weight[124][116],
reservoir_weight[124][117],
reservoir_weight[124][118],
reservoir_weight[124][119],
reservoir_weight[124][120],
reservoir_weight[124][121],
reservoir_weight[124][122],
reservoir_weight[124][123],
reservoir_weight[124][124],
reservoir_weight[124][125],
reservoir_weight[124][126],
reservoir_weight[124][127],
reservoir_weight[124][128],
reservoir_weight[124][129],
reservoir_weight[124][130],
reservoir_weight[124][131],
reservoir_weight[124][132],
reservoir_weight[124][133],
reservoir_weight[124][134],
reservoir_weight[124][135],
reservoir_weight[124][136],
reservoir_weight[124][137],
reservoir_weight[124][138],
reservoir_weight[124][139],
reservoir_weight[124][140],
reservoir_weight[124][141],
reservoir_weight[124][142],
reservoir_weight[124][143],
reservoir_weight[124][144],
reservoir_weight[124][145],
reservoir_weight[124][146],
reservoir_weight[124][147],
reservoir_weight[124][148],
reservoir_weight[124][149],
reservoir_weight[124][150],
reservoir_weight[124][151],
reservoir_weight[124][152],
reservoir_weight[124][153],
reservoir_weight[124][154],
reservoir_weight[124][155],
reservoir_weight[124][156],
reservoir_weight[124][157],
reservoir_weight[124][158],
reservoir_weight[124][159],
reservoir_weight[124][160],
reservoir_weight[124][161],
reservoir_weight[124][162],
reservoir_weight[124][163],
reservoir_weight[124][164],
reservoir_weight[124][165],
reservoir_weight[124][166],
reservoir_weight[124][167],
reservoir_weight[124][168],
reservoir_weight[124][169],
reservoir_weight[124][170],
reservoir_weight[124][171],
reservoir_weight[124][172],
reservoir_weight[124][173],
reservoir_weight[124][174],
reservoir_weight[124][175],
reservoir_weight[124][176],
reservoir_weight[124][177],
reservoir_weight[124][178],
reservoir_weight[124][179],
reservoir_weight[124][180],
reservoir_weight[124][181],
reservoir_weight[124][182],
reservoir_weight[124][183],
reservoir_weight[124][184],
reservoir_weight[124][185],
reservoir_weight[124][186],
reservoir_weight[124][187],
reservoir_weight[124][188],
reservoir_weight[124][189],
reservoir_weight[124][190],
reservoir_weight[124][191],
reservoir_weight[124][192],
reservoir_weight[124][193],
reservoir_weight[124][194],
reservoir_weight[124][195],
reservoir_weight[124][196],
reservoir_weight[124][197],
reservoir_weight[124][198],
reservoir_weight[124][199]
},
{reservoir_weight[125][0],
reservoir_weight[125][1],
reservoir_weight[125][2],
reservoir_weight[125][3],
reservoir_weight[125][4],
reservoir_weight[125][5],
reservoir_weight[125][6],
reservoir_weight[125][7],
reservoir_weight[125][8],
reservoir_weight[125][9],
reservoir_weight[125][10],
reservoir_weight[125][11],
reservoir_weight[125][12],
reservoir_weight[125][13],
reservoir_weight[125][14],
reservoir_weight[125][15],
reservoir_weight[125][16],
reservoir_weight[125][17],
reservoir_weight[125][18],
reservoir_weight[125][19],
reservoir_weight[125][20],
reservoir_weight[125][21],
reservoir_weight[125][22],
reservoir_weight[125][23],
reservoir_weight[125][24],
reservoir_weight[125][25],
reservoir_weight[125][26],
reservoir_weight[125][27],
reservoir_weight[125][28],
reservoir_weight[125][29],
reservoir_weight[125][30],
reservoir_weight[125][31],
reservoir_weight[125][32],
reservoir_weight[125][33],
reservoir_weight[125][34],
reservoir_weight[125][35],
reservoir_weight[125][36],
reservoir_weight[125][37],
reservoir_weight[125][38],
reservoir_weight[125][39],
reservoir_weight[125][40],
reservoir_weight[125][41],
reservoir_weight[125][42],
reservoir_weight[125][43],
reservoir_weight[125][44],
reservoir_weight[125][45],
reservoir_weight[125][46],
reservoir_weight[125][47],
reservoir_weight[125][48],
reservoir_weight[125][49],
reservoir_weight[125][50],
reservoir_weight[125][51],
reservoir_weight[125][52],
reservoir_weight[125][53],
reservoir_weight[125][54],
reservoir_weight[125][55],
reservoir_weight[125][56],
reservoir_weight[125][57],
reservoir_weight[125][58],
reservoir_weight[125][59],
reservoir_weight[125][60],
reservoir_weight[125][61],
reservoir_weight[125][62],
reservoir_weight[125][63],
reservoir_weight[125][64],
reservoir_weight[125][65],
reservoir_weight[125][66],
reservoir_weight[125][67],
reservoir_weight[125][68],
reservoir_weight[125][69],
reservoir_weight[125][70],
reservoir_weight[125][71],
reservoir_weight[125][72],
reservoir_weight[125][73],
reservoir_weight[125][74],
reservoir_weight[125][75],
reservoir_weight[125][76],
reservoir_weight[125][77],
reservoir_weight[125][78],
reservoir_weight[125][79],
reservoir_weight[125][80],
reservoir_weight[125][81],
reservoir_weight[125][82],
reservoir_weight[125][83],
reservoir_weight[125][84],
reservoir_weight[125][85],
reservoir_weight[125][86],
reservoir_weight[125][87],
reservoir_weight[125][88],
reservoir_weight[125][89],
reservoir_weight[125][90],
reservoir_weight[125][91],
reservoir_weight[125][92],
reservoir_weight[125][93],
reservoir_weight[125][94],
reservoir_weight[125][95],
reservoir_weight[125][96],
reservoir_weight[125][97],
reservoir_weight[125][98],
reservoir_weight[125][99],
reservoir_weight[125][100],
reservoir_weight[125][101],
reservoir_weight[125][102],
reservoir_weight[125][103],
reservoir_weight[125][104],
reservoir_weight[125][105],
reservoir_weight[125][106],
reservoir_weight[125][107],
reservoir_weight[125][108],
reservoir_weight[125][109],
reservoir_weight[125][110],
reservoir_weight[125][111],
reservoir_weight[125][112],
reservoir_weight[125][113],
reservoir_weight[125][114],
reservoir_weight[125][115],
reservoir_weight[125][116],
reservoir_weight[125][117],
reservoir_weight[125][118],
reservoir_weight[125][119],
reservoir_weight[125][120],
reservoir_weight[125][121],
reservoir_weight[125][122],
reservoir_weight[125][123],
reservoir_weight[125][124],
reservoir_weight[125][125],
reservoir_weight[125][126],
reservoir_weight[125][127],
reservoir_weight[125][128],
reservoir_weight[125][129],
reservoir_weight[125][130],
reservoir_weight[125][131],
reservoir_weight[125][132],
reservoir_weight[125][133],
reservoir_weight[125][134],
reservoir_weight[125][135],
reservoir_weight[125][136],
reservoir_weight[125][137],
reservoir_weight[125][138],
reservoir_weight[125][139],
reservoir_weight[125][140],
reservoir_weight[125][141],
reservoir_weight[125][142],
reservoir_weight[125][143],
reservoir_weight[125][144],
reservoir_weight[125][145],
reservoir_weight[125][146],
reservoir_weight[125][147],
reservoir_weight[125][148],
reservoir_weight[125][149],
reservoir_weight[125][150],
reservoir_weight[125][151],
reservoir_weight[125][152],
reservoir_weight[125][153],
reservoir_weight[125][154],
reservoir_weight[125][155],
reservoir_weight[125][156],
reservoir_weight[125][157],
reservoir_weight[125][158],
reservoir_weight[125][159],
reservoir_weight[125][160],
reservoir_weight[125][161],
reservoir_weight[125][162],
reservoir_weight[125][163],
reservoir_weight[125][164],
reservoir_weight[125][165],
reservoir_weight[125][166],
reservoir_weight[125][167],
reservoir_weight[125][168],
reservoir_weight[125][169],
reservoir_weight[125][170],
reservoir_weight[125][171],
reservoir_weight[125][172],
reservoir_weight[125][173],
reservoir_weight[125][174],
reservoir_weight[125][175],
reservoir_weight[125][176],
reservoir_weight[125][177],
reservoir_weight[125][178],
reservoir_weight[125][179],
reservoir_weight[125][180],
reservoir_weight[125][181],
reservoir_weight[125][182],
reservoir_weight[125][183],
reservoir_weight[125][184],
reservoir_weight[125][185],
reservoir_weight[125][186],
reservoir_weight[125][187],
reservoir_weight[125][188],
reservoir_weight[125][189],
reservoir_weight[125][190],
reservoir_weight[125][191],
reservoir_weight[125][192],
reservoir_weight[125][193],
reservoir_weight[125][194],
reservoir_weight[125][195],
reservoir_weight[125][196],
reservoir_weight[125][197],
reservoir_weight[125][198],
reservoir_weight[125][199]
},
{reservoir_weight[126][0],
reservoir_weight[126][1],
reservoir_weight[126][2],
reservoir_weight[126][3],
reservoir_weight[126][4],
reservoir_weight[126][5],
reservoir_weight[126][6],
reservoir_weight[126][7],
reservoir_weight[126][8],
reservoir_weight[126][9],
reservoir_weight[126][10],
reservoir_weight[126][11],
reservoir_weight[126][12],
reservoir_weight[126][13],
reservoir_weight[126][14],
reservoir_weight[126][15],
reservoir_weight[126][16],
reservoir_weight[126][17],
reservoir_weight[126][18],
reservoir_weight[126][19],
reservoir_weight[126][20],
reservoir_weight[126][21],
reservoir_weight[126][22],
reservoir_weight[126][23],
reservoir_weight[126][24],
reservoir_weight[126][25],
reservoir_weight[126][26],
reservoir_weight[126][27],
reservoir_weight[126][28],
reservoir_weight[126][29],
reservoir_weight[126][30],
reservoir_weight[126][31],
reservoir_weight[126][32],
reservoir_weight[126][33],
reservoir_weight[126][34],
reservoir_weight[126][35],
reservoir_weight[126][36],
reservoir_weight[126][37],
reservoir_weight[126][38],
reservoir_weight[126][39],
reservoir_weight[126][40],
reservoir_weight[126][41],
reservoir_weight[126][42],
reservoir_weight[126][43],
reservoir_weight[126][44],
reservoir_weight[126][45],
reservoir_weight[126][46],
reservoir_weight[126][47],
reservoir_weight[126][48],
reservoir_weight[126][49],
reservoir_weight[126][50],
reservoir_weight[126][51],
reservoir_weight[126][52],
reservoir_weight[126][53],
reservoir_weight[126][54],
reservoir_weight[126][55],
reservoir_weight[126][56],
reservoir_weight[126][57],
reservoir_weight[126][58],
reservoir_weight[126][59],
reservoir_weight[126][60],
reservoir_weight[126][61],
reservoir_weight[126][62],
reservoir_weight[126][63],
reservoir_weight[126][64],
reservoir_weight[126][65],
reservoir_weight[126][66],
reservoir_weight[126][67],
reservoir_weight[126][68],
reservoir_weight[126][69],
reservoir_weight[126][70],
reservoir_weight[126][71],
reservoir_weight[126][72],
reservoir_weight[126][73],
reservoir_weight[126][74],
reservoir_weight[126][75],
reservoir_weight[126][76],
reservoir_weight[126][77],
reservoir_weight[126][78],
reservoir_weight[126][79],
reservoir_weight[126][80],
reservoir_weight[126][81],
reservoir_weight[126][82],
reservoir_weight[126][83],
reservoir_weight[126][84],
reservoir_weight[126][85],
reservoir_weight[126][86],
reservoir_weight[126][87],
reservoir_weight[126][88],
reservoir_weight[126][89],
reservoir_weight[126][90],
reservoir_weight[126][91],
reservoir_weight[126][92],
reservoir_weight[126][93],
reservoir_weight[126][94],
reservoir_weight[126][95],
reservoir_weight[126][96],
reservoir_weight[126][97],
reservoir_weight[126][98],
reservoir_weight[126][99],
reservoir_weight[126][100],
reservoir_weight[126][101],
reservoir_weight[126][102],
reservoir_weight[126][103],
reservoir_weight[126][104],
reservoir_weight[126][105],
reservoir_weight[126][106],
reservoir_weight[126][107],
reservoir_weight[126][108],
reservoir_weight[126][109],
reservoir_weight[126][110],
reservoir_weight[126][111],
reservoir_weight[126][112],
reservoir_weight[126][113],
reservoir_weight[126][114],
reservoir_weight[126][115],
reservoir_weight[126][116],
reservoir_weight[126][117],
reservoir_weight[126][118],
reservoir_weight[126][119],
reservoir_weight[126][120],
reservoir_weight[126][121],
reservoir_weight[126][122],
reservoir_weight[126][123],
reservoir_weight[126][124],
reservoir_weight[126][125],
reservoir_weight[126][126],
reservoir_weight[126][127],
reservoir_weight[126][128],
reservoir_weight[126][129],
reservoir_weight[126][130],
reservoir_weight[126][131],
reservoir_weight[126][132],
reservoir_weight[126][133],
reservoir_weight[126][134],
reservoir_weight[126][135],
reservoir_weight[126][136],
reservoir_weight[126][137],
reservoir_weight[126][138],
reservoir_weight[126][139],
reservoir_weight[126][140],
reservoir_weight[126][141],
reservoir_weight[126][142],
reservoir_weight[126][143],
reservoir_weight[126][144],
reservoir_weight[126][145],
reservoir_weight[126][146],
reservoir_weight[126][147],
reservoir_weight[126][148],
reservoir_weight[126][149],
reservoir_weight[126][150],
reservoir_weight[126][151],
reservoir_weight[126][152],
reservoir_weight[126][153],
reservoir_weight[126][154],
reservoir_weight[126][155],
reservoir_weight[126][156],
reservoir_weight[126][157],
reservoir_weight[126][158],
reservoir_weight[126][159],
reservoir_weight[126][160],
reservoir_weight[126][161],
reservoir_weight[126][162],
reservoir_weight[126][163],
reservoir_weight[126][164],
reservoir_weight[126][165],
reservoir_weight[126][166],
reservoir_weight[126][167],
reservoir_weight[126][168],
reservoir_weight[126][169],
reservoir_weight[126][170],
reservoir_weight[126][171],
reservoir_weight[126][172],
reservoir_weight[126][173],
reservoir_weight[126][174],
reservoir_weight[126][175],
reservoir_weight[126][176],
reservoir_weight[126][177],
reservoir_weight[126][178],
reservoir_weight[126][179],
reservoir_weight[126][180],
reservoir_weight[126][181],
reservoir_weight[126][182],
reservoir_weight[126][183],
reservoir_weight[126][184],
reservoir_weight[126][185],
reservoir_weight[126][186],
reservoir_weight[126][187],
reservoir_weight[126][188],
reservoir_weight[126][189],
reservoir_weight[126][190],
reservoir_weight[126][191],
reservoir_weight[126][192],
reservoir_weight[126][193],
reservoir_weight[126][194],
reservoir_weight[126][195],
reservoir_weight[126][196],
reservoir_weight[126][197],
reservoir_weight[126][198],
reservoir_weight[126][199]
},
{reservoir_weight[127][0],
reservoir_weight[127][1],
reservoir_weight[127][2],
reservoir_weight[127][3],
reservoir_weight[127][4],
reservoir_weight[127][5],
reservoir_weight[127][6],
reservoir_weight[127][7],
reservoir_weight[127][8],
reservoir_weight[127][9],
reservoir_weight[127][10],
reservoir_weight[127][11],
reservoir_weight[127][12],
reservoir_weight[127][13],
reservoir_weight[127][14],
reservoir_weight[127][15],
reservoir_weight[127][16],
reservoir_weight[127][17],
reservoir_weight[127][18],
reservoir_weight[127][19],
reservoir_weight[127][20],
reservoir_weight[127][21],
reservoir_weight[127][22],
reservoir_weight[127][23],
reservoir_weight[127][24],
reservoir_weight[127][25],
reservoir_weight[127][26],
reservoir_weight[127][27],
reservoir_weight[127][28],
reservoir_weight[127][29],
reservoir_weight[127][30],
reservoir_weight[127][31],
reservoir_weight[127][32],
reservoir_weight[127][33],
reservoir_weight[127][34],
reservoir_weight[127][35],
reservoir_weight[127][36],
reservoir_weight[127][37],
reservoir_weight[127][38],
reservoir_weight[127][39],
reservoir_weight[127][40],
reservoir_weight[127][41],
reservoir_weight[127][42],
reservoir_weight[127][43],
reservoir_weight[127][44],
reservoir_weight[127][45],
reservoir_weight[127][46],
reservoir_weight[127][47],
reservoir_weight[127][48],
reservoir_weight[127][49],
reservoir_weight[127][50],
reservoir_weight[127][51],
reservoir_weight[127][52],
reservoir_weight[127][53],
reservoir_weight[127][54],
reservoir_weight[127][55],
reservoir_weight[127][56],
reservoir_weight[127][57],
reservoir_weight[127][58],
reservoir_weight[127][59],
reservoir_weight[127][60],
reservoir_weight[127][61],
reservoir_weight[127][62],
reservoir_weight[127][63],
reservoir_weight[127][64],
reservoir_weight[127][65],
reservoir_weight[127][66],
reservoir_weight[127][67],
reservoir_weight[127][68],
reservoir_weight[127][69],
reservoir_weight[127][70],
reservoir_weight[127][71],
reservoir_weight[127][72],
reservoir_weight[127][73],
reservoir_weight[127][74],
reservoir_weight[127][75],
reservoir_weight[127][76],
reservoir_weight[127][77],
reservoir_weight[127][78],
reservoir_weight[127][79],
reservoir_weight[127][80],
reservoir_weight[127][81],
reservoir_weight[127][82],
reservoir_weight[127][83],
reservoir_weight[127][84],
reservoir_weight[127][85],
reservoir_weight[127][86],
reservoir_weight[127][87],
reservoir_weight[127][88],
reservoir_weight[127][89],
reservoir_weight[127][90],
reservoir_weight[127][91],
reservoir_weight[127][92],
reservoir_weight[127][93],
reservoir_weight[127][94],
reservoir_weight[127][95],
reservoir_weight[127][96],
reservoir_weight[127][97],
reservoir_weight[127][98],
reservoir_weight[127][99],
reservoir_weight[127][100],
reservoir_weight[127][101],
reservoir_weight[127][102],
reservoir_weight[127][103],
reservoir_weight[127][104],
reservoir_weight[127][105],
reservoir_weight[127][106],
reservoir_weight[127][107],
reservoir_weight[127][108],
reservoir_weight[127][109],
reservoir_weight[127][110],
reservoir_weight[127][111],
reservoir_weight[127][112],
reservoir_weight[127][113],
reservoir_weight[127][114],
reservoir_weight[127][115],
reservoir_weight[127][116],
reservoir_weight[127][117],
reservoir_weight[127][118],
reservoir_weight[127][119],
reservoir_weight[127][120],
reservoir_weight[127][121],
reservoir_weight[127][122],
reservoir_weight[127][123],
reservoir_weight[127][124],
reservoir_weight[127][125],
reservoir_weight[127][126],
reservoir_weight[127][127],
reservoir_weight[127][128],
reservoir_weight[127][129],
reservoir_weight[127][130],
reservoir_weight[127][131],
reservoir_weight[127][132],
reservoir_weight[127][133],
reservoir_weight[127][134],
reservoir_weight[127][135],
reservoir_weight[127][136],
reservoir_weight[127][137],
reservoir_weight[127][138],
reservoir_weight[127][139],
reservoir_weight[127][140],
reservoir_weight[127][141],
reservoir_weight[127][142],
reservoir_weight[127][143],
reservoir_weight[127][144],
reservoir_weight[127][145],
reservoir_weight[127][146],
reservoir_weight[127][147],
reservoir_weight[127][148],
reservoir_weight[127][149],
reservoir_weight[127][150],
reservoir_weight[127][151],
reservoir_weight[127][152],
reservoir_weight[127][153],
reservoir_weight[127][154],
reservoir_weight[127][155],
reservoir_weight[127][156],
reservoir_weight[127][157],
reservoir_weight[127][158],
reservoir_weight[127][159],
reservoir_weight[127][160],
reservoir_weight[127][161],
reservoir_weight[127][162],
reservoir_weight[127][163],
reservoir_weight[127][164],
reservoir_weight[127][165],
reservoir_weight[127][166],
reservoir_weight[127][167],
reservoir_weight[127][168],
reservoir_weight[127][169],
reservoir_weight[127][170],
reservoir_weight[127][171],
reservoir_weight[127][172],
reservoir_weight[127][173],
reservoir_weight[127][174],
reservoir_weight[127][175],
reservoir_weight[127][176],
reservoir_weight[127][177],
reservoir_weight[127][178],
reservoir_weight[127][179],
reservoir_weight[127][180],
reservoir_weight[127][181],
reservoir_weight[127][182],
reservoir_weight[127][183],
reservoir_weight[127][184],
reservoir_weight[127][185],
reservoir_weight[127][186],
reservoir_weight[127][187],
reservoir_weight[127][188],
reservoir_weight[127][189],
reservoir_weight[127][190],
reservoir_weight[127][191],
reservoir_weight[127][192],
reservoir_weight[127][193],
reservoir_weight[127][194],
reservoir_weight[127][195],
reservoir_weight[127][196],
reservoir_weight[127][197],
reservoir_weight[127][198],
reservoir_weight[127][199]
},
{reservoir_weight[128][0],
reservoir_weight[128][1],
reservoir_weight[128][2],
reservoir_weight[128][3],
reservoir_weight[128][4],
reservoir_weight[128][5],
reservoir_weight[128][6],
reservoir_weight[128][7],
reservoir_weight[128][8],
reservoir_weight[128][9],
reservoir_weight[128][10],
reservoir_weight[128][11],
reservoir_weight[128][12],
reservoir_weight[128][13],
reservoir_weight[128][14],
reservoir_weight[128][15],
reservoir_weight[128][16],
reservoir_weight[128][17],
reservoir_weight[128][18],
reservoir_weight[128][19],
reservoir_weight[128][20],
reservoir_weight[128][21],
reservoir_weight[128][22],
reservoir_weight[128][23],
reservoir_weight[128][24],
reservoir_weight[128][25],
reservoir_weight[128][26],
reservoir_weight[128][27],
reservoir_weight[128][28],
reservoir_weight[128][29],
reservoir_weight[128][30],
reservoir_weight[128][31],
reservoir_weight[128][32],
reservoir_weight[128][33],
reservoir_weight[128][34],
reservoir_weight[128][35],
reservoir_weight[128][36],
reservoir_weight[128][37],
reservoir_weight[128][38],
reservoir_weight[128][39],
reservoir_weight[128][40],
reservoir_weight[128][41],
reservoir_weight[128][42],
reservoir_weight[128][43],
reservoir_weight[128][44],
reservoir_weight[128][45],
reservoir_weight[128][46],
reservoir_weight[128][47],
reservoir_weight[128][48],
reservoir_weight[128][49],
reservoir_weight[128][50],
reservoir_weight[128][51],
reservoir_weight[128][52],
reservoir_weight[128][53],
reservoir_weight[128][54],
reservoir_weight[128][55],
reservoir_weight[128][56],
reservoir_weight[128][57],
reservoir_weight[128][58],
reservoir_weight[128][59],
reservoir_weight[128][60],
reservoir_weight[128][61],
reservoir_weight[128][62],
reservoir_weight[128][63],
reservoir_weight[128][64],
reservoir_weight[128][65],
reservoir_weight[128][66],
reservoir_weight[128][67],
reservoir_weight[128][68],
reservoir_weight[128][69],
reservoir_weight[128][70],
reservoir_weight[128][71],
reservoir_weight[128][72],
reservoir_weight[128][73],
reservoir_weight[128][74],
reservoir_weight[128][75],
reservoir_weight[128][76],
reservoir_weight[128][77],
reservoir_weight[128][78],
reservoir_weight[128][79],
reservoir_weight[128][80],
reservoir_weight[128][81],
reservoir_weight[128][82],
reservoir_weight[128][83],
reservoir_weight[128][84],
reservoir_weight[128][85],
reservoir_weight[128][86],
reservoir_weight[128][87],
reservoir_weight[128][88],
reservoir_weight[128][89],
reservoir_weight[128][90],
reservoir_weight[128][91],
reservoir_weight[128][92],
reservoir_weight[128][93],
reservoir_weight[128][94],
reservoir_weight[128][95],
reservoir_weight[128][96],
reservoir_weight[128][97],
reservoir_weight[128][98],
reservoir_weight[128][99],
reservoir_weight[128][100],
reservoir_weight[128][101],
reservoir_weight[128][102],
reservoir_weight[128][103],
reservoir_weight[128][104],
reservoir_weight[128][105],
reservoir_weight[128][106],
reservoir_weight[128][107],
reservoir_weight[128][108],
reservoir_weight[128][109],
reservoir_weight[128][110],
reservoir_weight[128][111],
reservoir_weight[128][112],
reservoir_weight[128][113],
reservoir_weight[128][114],
reservoir_weight[128][115],
reservoir_weight[128][116],
reservoir_weight[128][117],
reservoir_weight[128][118],
reservoir_weight[128][119],
reservoir_weight[128][120],
reservoir_weight[128][121],
reservoir_weight[128][122],
reservoir_weight[128][123],
reservoir_weight[128][124],
reservoir_weight[128][125],
reservoir_weight[128][126],
reservoir_weight[128][127],
reservoir_weight[128][128],
reservoir_weight[128][129],
reservoir_weight[128][130],
reservoir_weight[128][131],
reservoir_weight[128][132],
reservoir_weight[128][133],
reservoir_weight[128][134],
reservoir_weight[128][135],
reservoir_weight[128][136],
reservoir_weight[128][137],
reservoir_weight[128][138],
reservoir_weight[128][139],
reservoir_weight[128][140],
reservoir_weight[128][141],
reservoir_weight[128][142],
reservoir_weight[128][143],
reservoir_weight[128][144],
reservoir_weight[128][145],
reservoir_weight[128][146],
reservoir_weight[128][147],
reservoir_weight[128][148],
reservoir_weight[128][149],
reservoir_weight[128][150],
reservoir_weight[128][151],
reservoir_weight[128][152],
reservoir_weight[128][153],
reservoir_weight[128][154],
reservoir_weight[128][155],
reservoir_weight[128][156],
reservoir_weight[128][157],
reservoir_weight[128][158],
reservoir_weight[128][159],
reservoir_weight[128][160],
reservoir_weight[128][161],
reservoir_weight[128][162],
reservoir_weight[128][163],
reservoir_weight[128][164],
reservoir_weight[128][165],
reservoir_weight[128][166],
reservoir_weight[128][167],
reservoir_weight[128][168],
reservoir_weight[128][169],
reservoir_weight[128][170],
reservoir_weight[128][171],
reservoir_weight[128][172],
reservoir_weight[128][173],
reservoir_weight[128][174],
reservoir_weight[128][175],
reservoir_weight[128][176],
reservoir_weight[128][177],
reservoir_weight[128][178],
reservoir_weight[128][179],
reservoir_weight[128][180],
reservoir_weight[128][181],
reservoir_weight[128][182],
reservoir_weight[128][183],
reservoir_weight[128][184],
reservoir_weight[128][185],
reservoir_weight[128][186],
reservoir_weight[128][187],
reservoir_weight[128][188],
reservoir_weight[128][189],
reservoir_weight[128][190],
reservoir_weight[128][191],
reservoir_weight[128][192],
reservoir_weight[128][193],
reservoir_weight[128][194],
reservoir_weight[128][195],
reservoir_weight[128][196],
reservoir_weight[128][197],
reservoir_weight[128][198],
reservoir_weight[128][199]
},
{reservoir_weight[129][0],
reservoir_weight[129][1],
reservoir_weight[129][2],
reservoir_weight[129][3],
reservoir_weight[129][4],
reservoir_weight[129][5],
reservoir_weight[129][6],
reservoir_weight[129][7],
reservoir_weight[129][8],
reservoir_weight[129][9],
reservoir_weight[129][10],
reservoir_weight[129][11],
reservoir_weight[129][12],
reservoir_weight[129][13],
reservoir_weight[129][14],
reservoir_weight[129][15],
reservoir_weight[129][16],
reservoir_weight[129][17],
reservoir_weight[129][18],
reservoir_weight[129][19],
reservoir_weight[129][20],
reservoir_weight[129][21],
reservoir_weight[129][22],
reservoir_weight[129][23],
reservoir_weight[129][24],
reservoir_weight[129][25],
reservoir_weight[129][26],
reservoir_weight[129][27],
reservoir_weight[129][28],
reservoir_weight[129][29],
reservoir_weight[129][30],
reservoir_weight[129][31],
reservoir_weight[129][32],
reservoir_weight[129][33],
reservoir_weight[129][34],
reservoir_weight[129][35],
reservoir_weight[129][36],
reservoir_weight[129][37],
reservoir_weight[129][38],
reservoir_weight[129][39],
reservoir_weight[129][40],
reservoir_weight[129][41],
reservoir_weight[129][42],
reservoir_weight[129][43],
reservoir_weight[129][44],
reservoir_weight[129][45],
reservoir_weight[129][46],
reservoir_weight[129][47],
reservoir_weight[129][48],
reservoir_weight[129][49],
reservoir_weight[129][50],
reservoir_weight[129][51],
reservoir_weight[129][52],
reservoir_weight[129][53],
reservoir_weight[129][54],
reservoir_weight[129][55],
reservoir_weight[129][56],
reservoir_weight[129][57],
reservoir_weight[129][58],
reservoir_weight[129][59],
reservoir_weight[129][60],
reservoir_weight[129][61],
reservoir_weight[129][62],
reservoir_weight[129][63],
reservoir_weight[129][64],
reservoir_weight[129][65],
reservoir_weight[129][66],
reservoir_weight[129][67],
reservoir_weight[129][68],
reservoir_weight[129][69],
reservoir_weight[129][70],
reservoir_weight[129][71],
reservoir_weight[129][72],
reservoir_weight[129][73],
reservoir_weight[129][74],
reservoir_weight[129][75],
reservoir_weight[129][76],
reservoir_weight[129][77],
reservoir_weight[129][78],
reservoir_weight[129][79],
reservoir_weight[129][80],
reservoir_weight[129][81],
reservoir_weight[129][82],
reservoir_weight[129][83],
reservoir_weight[129][84],
reservoir_weight[129][85],
reservoir_weight[129][86],
reservoir_weight[129][87],
reservoir_weight[129][88],
reservoir_weight[129][89],
reservoir_weight[129][90],
reservoir_weight[129][91],
reservoir_weight[129][92],
reservoir_weight[129][93],
reservoir_weight[129][94],
reservoir_weight[129][95],
reservoir_weight[129][96],
reservoir_weight[129][97],
reservoir_weight[129][98],
reservoir_weight[129][99],
reservoir_weight[129][100],
reservoir_weight[129][101],
reservoir_weight[129][102],
reservoir_weight[129][103],
reservoir_weight[129][104],
reservoir_weight[129][105],
reservoir_weight[129][106],
reservoir_weight[129][107],
reservoir_weight[129][108],
reservoir_weight[129][109],
reservoir_weight[129][110],
reservoir_weight[129][111],
reservoir_weight[129][112],
reservoir_weight[129][113],
reservoir_weight[129][114],
reservoir_weight[129][115],
reservoir_weight[129][116],
reservoir_weight[129][117],
reservoir_weight[129][118],
reservoir_weight[129][119],
reservoir_weight[129][120],
reservoir_weight[129][121],
reservoir_weight[129][122],
reservoir_weight[129][123],
reservoir_weight[129][124],
reservoir_weight[129][125],
reservoir_weight[129][126],
reservoir_weight[129][127],
reservoir_weight[129][128],
reservoir_weight[129][129],
reservoir_weight[129][130],
reservoir_weight[129][131],
reservoir_weight[129][132],
reservoir_weight[129][133],
reservoir_weight[129][134],
reservoir_weight[129][135],
reservoir_weight[129][136],
reservoir_weight[129][137],
reservoir_weight[129][138],
reservoir_weight[129][139],
reservoir_weight[129][140],
reservoir_weight[129][141],
reservoir_weight[129][142],
reservoir_weight[129][143],
reservoir_weight[129][144],
reservoir_weight[129][145],
reservoir_weight[129][146],
reservoir_weight[129][147],
reservoir_weight[129][148],
reservoir_weight[129][149],
reservoir_weight[129][150],
reservoir_weight[129][151],
reservoir_weight[129][152],
reservoir_weight[129][153],
reservoir_weight[129][154],
reservoir_weight[129][155],
reservoir_weight[129][156],
reservoir_weight[129][157],
reservoir_weight[129][158],
reservoir_weight[129][159],
reservoir_weight[129][160],
reservoir_weight[129][161],
reservoir_weight[129][162],
reservoir_weight[129][163],
reservoir_weight[129][164],
reservoir_weight[129][165],
reservoir_weight[129][166],
reservoir_weight[129][167],
reservoir_weight[129][168],
reservoir_weight[129][169],
reservoir_weight[129][170],
reservoir_weight[129][171],
reservoir_weight[129][172],
reservoir_weight[129][173],
reservoir_weight[129][174],
reservoir_weight[129][175],
reservoir_weight[129][176],
reservoir_weight[129][177],
reservoir_weight[129][178],
reservoir_weight[129][179],
reservoir_weight[129][180],
reservoir_weight[129][181],
reservoir_weight[129][182],
reservoir_weight[129][183],
reservoir_weight[129][184],
reservoir_weight[129][185],
reservoir_weight[129][186],
reservoir_weight[129][187],
reservoir_weight[129][188],
reservoir_weight[129][189],
reservoir_weight[129][190],
reservoir_weight[129][191],
reservoir_weight[129][192],
reservoir_weight[129][193],
reservoir_weight[129][194],
reservoir_weight[129][195],
reservoir_weight[129][196],
reservoir_weight[129][197],
reservoir_weight[129][198],
reservoir_weight[129][199]
},
{reservoir_weight[130][0],
reservoir_weight[130][1],
reservoir_weight[130][2],
reservoir_weight[130][3],
reservoir_weight[130][4],
reservoir_weight[130][5],
reservoir_weight[130][6],
reservoir_weight[130][7],
reservoir_weight[130][8],
reservoir_weight[130][9],
reservoir_weight[130][10],
reservoir_weight[130][11],
reservoir_weight[130][12],
reservoir_weight[130][13],
reservoir_weight[130][14],
reservoir_weight[130][15],
reservoir_weight[130][16],
reservoir_weight[130][17],
reservoir_weight[130][18],
reservoir_weight[130][19],
reservoir_weight[130][20],
reservoir_weight[130][21],
reservoir_weight[130][22],
reservoir_weight[130][23],
reservoir_weight[130][24],
reservoir_weight[130][25],
reservoir_weight[130][26],
reservoir_weight[130][27],
reservoir_weight[130][28],
reservoir_weight[130][29],
reservoir_weight[130][30],
reservoir_weight[130][31],
reservoir_weight[130][32],
reservoir_weight[130][33],
reservoir_weight[130][34],
reservoir_weight[130][35],
reservoir_weight[130][36],
reservoir_weight[130][37],
reservoir_weight[130][38],
reservoir_weight[130][39],
reservoir_weight[130][40],
reservoir_weight[130][41],
reservoir_weight[130][42],
reservoir_weight[130][43],
reservoir_weight[130][44],
reservoir_weight[130][45],
reservoir_weight[130][46],
reservoir_weight[130][47],
reservoir_weight[130][48],
reservoir_weight[130][49],
reservoir_weight[130][50],
reservoir_weight[130][51],
reservoir_weight[130][52],
reservoir_weight[130][53],
reservoir_weight[130][54],
reservoir_weight[130][55],
reservoir_weight[130][56],
reservoir_weight[130][57],
reservoir_weight[130][58],
reservoir_weight[130][59],
reservoir_weight[130][60],
reservoir_weight[130][61],
reservoir_weight[130][62],
reservoir_weight[130][63],
reservoir_weight[130][64],
reservoir_weight[130][65],
reservoir_weight[130][66],
reservoir_weight[130][67],
reservoir_weight[130][68],
reservoir_weight[130][69],
reservoir_weight[130][70],
reservoir_weight[130][71],
reservoir_weight[130][72],
reservoir_weight[130][73],
reservoir_weight[130][74],
reservoir_weight[130][75],
reservoir_weight[130][76],
reservoir_weight[130][77],
reservoir_weight[130][78],
reservoir_weight[130][79],
reservoir_weight[130][80],
reservoir_weight[130][81],
reservoir_weight[130][82],
reservoir_weight[130][83],
reservoir_weight[130][84],
reservoir_weight[130][85],
reservoir_weight[130][86],
reservoir_weight[130][87],
reservoir_weight[130][88],
reservoir_weight[130][89],
reservoir_weight[130][90],
reservoir_weight[130][91],
reservoir_weight[130][92],
reservoir_weight[130][93],
reservoir_weight[130][94],
reservoir_weight[130][95],
reservoir_weight[130][96],
reservoir_weight[130][97],
reservoir_weight[130][98],
reservoir_weight[130][99],
reservoir_weight[130][100],
reservoir_weight[130][101],
reservoir_weight[130][102],
reservoir_weight[130][103],
reservoir_weight[130][104],
reservoir_weight[130][105],
reservoir_weight[130][106],
reservoir_weight[130][107],
reservoir_weight[130][108],
reservoir_weight[130][109],
reservoir_weight[130][110],
reservoir_weight[130][111],
reservoir_weight[130][112],
reservoir_weight[130][113],
reservoir_weight[130][114],
reservoir_weight[130][115],
reservoir_weight[130][116],
reservoir_weight[130][117],
reservoir_weight[130][118],
reservoir_weight[130][119],
reservoir_weight[130][120],
reservoir_weight[130][121],
reservoir_weight[130][122],
reservoir_weight[130][123],
reservoir_weight[130][124],
reservoir_weight[130][125],
reservoir_weight[130][126],
reservoir_weight[130][127],
reservoir_weight[130][128],
reservoir_weight[130][129],
reservoir_weight[130][130],
reservoir_weight[130][131],
reservoir_weight[130][132],
reservoir_weight[130][133],
reservoir_weight[130][134],
reservoir_weight[130][135],
reservoir_weight[130][136],
reservoir_weight[130][137],
reservoir_weight[130][138],
reservoir_weight[130][139],
reservoir_weight[130][140],
reservoir_weight[130][141],
reservoir_weight[130][142],
reservoir_weight[130][143],
reservoir_weight[130][144],
reservoir_weight[130][145],
reservoir_weight[130][146],
reservoir_weight[130][147],
reservoir_weight[130][148],
reservoir_weight[130][149],
reservoir_weight[130][150],
reservoir_weight[130][151],
reservoir_weight[130][152],
reservoir_weight[130][153],
reservoir_weight[130][154],
reservoir_weight[130][155],
reservoir_weight[130][156],
reservoir_weight[130][157],
reservoir_weight[130][158],
reservoir_weight[130][159],
reservoir_weight[130][160],
reservoir_weight[130][161],
reservoir_weight[130][162],
reservoir_weight[130][163],
reservoir_weight[130][164],
reservoir_weight[130][165],
reservoir_weight[130][166],
reservoir_weight[130][167],
reservoir_weight[130][168],
reservoir_weight[130][169],
reservoir_weight[130][170],
reservoir_weight[130][171],
reservoir_weight[130][172],
reservoir_weight[130][173],
reservoir_weight[130][174],
reservoir_weight[130][175],
reservoir_weight[130][176],
reservoir_weight[130][177],
reservoir_weight[130][178],
reservoir_weight[130][179],
reservoir_weight[130][180],
reservoir_weight[130][181],
reservoir_weight[130][182],
reservoir_weight[130][183],
reservoir_weight[130][184],
reservoir_weight[130][185],
reservoir_weight[130][186],
reservoir_weight[130][187],
reservoir_weight[130][188],
reservoir_weight[130][189],
reservoir_weight[130][190],
reservoir_weight[130][191],
reservoir_weight[130][192],
reservoir_weight[130][193],
reservoir_weight[130][194],
reservoir_weight[130][195],
reservoir_weight[130][196],
reservoir_weight[130][197],
reservoir_weight[130][198],
reservoir_weight[130][199]
},
{reservoir_weight[131][0],
reservoir_weight[131][1],
reservoir_weight[131][2],
reservoir_weight[131][3],
reservoir_weight[131][4],
reservoir_weight[131][5],
reservoir_weight[131][6],
reservoir_weight[131][7],
reservoir_weight[131][8],
reservoir_weight[131][9],
reservoir_weight[131][10],
reservoir_weight[131][11],
reservoir_weight[131][12],
reservoir_weight[131][13],
reservoir_weight[131][14],
reservoir_weight[131][15],
reservoir_weight[131][16],
reservoir_weight[131][17],
reservoir_weight[131][18],
reservoir_weight[131][19],
reservoir_weight[131][20],
reservoir_weight[131][21],
reservoir_weight[131][22],
reservoir_weight[131][23],
reservoir_weight[131][24],
reservoir_weight[131][25],
reservoir_weight[131][26],
reservoir_weight[131][27],
reservoir_weight[131][28],
reservoir_weight[131][29],
reservoir_weight[131][30],
reservoir_weight[131][31],
reservoir_weight[131][32],
reservoir_weight[131][33],
reservoir_weight[131][34],
reservoir_weight[131][35],
reservoir_weight[131][36],
reservoir_weight[131][37],
reservoir_weight[131][38],
reservoir_weight[131][39],
reservoir_weight[131][40],
reservoir_weight[131][41],
reservoir_weight[131][42],
reservoir_weight[131][43],
reservoir_weight[131][44],
reservoir_weight[131][45],
reservoir_weight[131][46],
reservoir_weight[131][47],
reservoir_weight[131][48],
reservoir_weight[131][49],
reservoir_weight[131][50],
reservoir_weight[131][51],
reservoir_weight[131][52],
reservoir_weight[131][53],
reservoir_weight[131][54],
reservoir_weight[131][55],
reservoir_weight[131][56],
reservoir_weight[131][57],
reservoir_weight[131][58],
reservoir_weight[131][59],
reservoir_weight[131][60],
reservoir_weight[131][61],
reservoir_weight[131][62],
reservoir_weight[131][63],
reservoir_weight[131][64],
reservoir_weight[131][65],
reservoir_weight[131][66],
reservoir_weight[131][67],
reservoir_weight[131][68],
reservoir_weight[131][69],
reservoir_weight[131][70],
reservoir_weight[131][71],
reservoir_weight[131][72],
reservoir_weight[131][73],
reservoir_weight[131][74],
reservoir_weight[131][75],
reservoir_weight[131][76],
reservoir_weight[131][77],
reservoir_weight[131][78],
reservoir_weight[131][79],
reservoir_weight[131][80],
reservoir_weight[131][81],
reservoir_weight[131][82],
reservoir_weight[131][83],
reservoir_weight[131][84],
reservoir_weight[131][85],
reservoir_weight[131][86],
reservoir_weight[131][87],
reservoir_weight[131][88],
reservoir_weight[131][89],
reservoir_weight[131][90],
reservoir_weight[131][91],
reservoir_weight[131][92],
reservoir_weight[131][93],
reservoir_weight[131][94],
reservoir_weight[131][95],
reservoir_weight[131][96],
reservoir_weight[131][97],
reservoir_weight[131][98],
reservoir_weight[131][99],
reservoir_weight[131][100],
reservoir_weight[131][101],
reservoir_weight[131][102],
reservoir_weight[131][103],
reservoir_weight[131][104],
reservoir_weight[131][105],
reservoir_weight[131][106],
reservoir_weight[131][107],
reservoir_weight[131][108],
reservoir_weight[131][109],
reservoir_weight[131][110],
reservoir_weight[131][111],
reservoir_weight[131][112],
reservoir_weight[131][113],
reservoir_weight[131][114],
reservoir_weight[131][115],
reservoir_weight[131][116],
reservoir_weight[131][117],
reservoir_weight[131][118],
reservoir_weight[131][119],
reservoir_weight[131][120],
reservoir_weight[131][121],
reservoir_weight[131][122],
reservoir_weight[131][123],
reservoir_weight[131][124],
reservoir_weight[131][125],
reservoir_weight[131][126],
reservoir_weight[131][127],
reservoir_weight[131][128],
reservoir_weight[131][129],
reservoir_weight[131][130],
reservoir_weight[131][131],
reservoir_weight[131][132],
reservoir_weight[131][133],
reservoir_weight[131][134],
reservoir_weight[131][135],
reservoir_weight[131][136],
reservoir_weight[131][137],
reservoir_weight[131][138],
reservoir_weight[131][139],
reservoir_weight[131][140],
reservoir_weight[131][141],
reservoir_weight[131][142],
reservoir_weight[131][143],
reservoir_weight[131][144],
reservoir_weight[131][145],
reservoir_weight[131][146],
reservoir_weight[131][147],
reservoir_weight[131][148],
reservoir_weight[131][149],
reservoir_weight[131][150],
reservoir_weight[131][151],
reservoir_weight[131][152],
reservoir_weight[131][153],
reservoir_weight[131][154],
reservoir_weight[131][155],
reservoir_weight[131][156],
reservoir_weight[131][157],
reservoir_weight[131][158],
reservoir_weight[131][159],
reservoir_weight[131][160],
reservoir_weight[131][161],
reservoir_weight[131][162],
reservoir_weight[131][163],
reservoir_weight[131][164],
reservoir_weight[131][165],
reservoir_weight[131][166],
reservoir_weight[131][167],
reservoir_weight[131][168],
reservoir_weight[131][169],
reservoir_weight[131][170],
reservoir_weight[131][171],
reservoir_weight[131][172],
reservoir_weight[131][173],
reservoir_weight[131][174],
reservoir_weight[131][175],
reservoir_weight[131][176],
reservoir_weight[131][177],
reservoir_weight[131][178],
reservoir_weight[131][179],
reservoir_weight[131][180],
reservoir_weight[131][181],
reservoir_weight[131][182],
reservoir_weight[131][183],
reservoir_weight[131][184],
reservoir_weight[131][185],
reservoir_weight[131][186],
reservoir_weight[131][187],
reservoir_weight[131][188],
reservoir_weight[131][189],
reservoir_weight[131][190],
reservoir_weight[131][191],
reservoir_weight[131][192],
reservoir_weight[131][193],
reservoir_weight[131][194],
reservoir_weight[131][195],
reservoir_weight[131][196],
reservoir_weight[131][197],
reservoir_weight[131][198],
reservoir_weight[131][199]
},
{reservoir_weight[132][0],
reservoir_weight[132][1],
reservoir_weight[132][2],
reservoir_weight[132][3],
reservoir_weight[132][4],
reservoir_weight[132][5],
reservoir_weight[132][6],
reservoir_weight[132][7],
reservoir_weight[132][8],
reservoir_weight[132][9],
reservoir_weight[132][10],
reservoir_weight[132][11],
reservoir_weight[132][12],
reservoir_weight[132][13],
reservoir_weight[132][14],
reservoir_weight[132][15],
reservoir_weight[132][16],
reservoir_weight[132][17],
reservoir_weight[132][18],
reservoir_weight[132][19],
reservoir_weight[132][20],
reservoir_weight[132][21],
reservoir_weight[132][22],
reservoir_weight[132][23],
reservoir_weight[132][24],
reservoir_weight[132][25],
reservoir_weight[132][26],
reservoir_weight[132][27],
reservoir_weight[132][28],
reservoir_weight[132][29],
reservoir_weight[132][30],
reservoir_weight[132][31],
reservoir_weight[132][32],
reservoir_weight[132][33],
reservoir_weight[132][34],
reservoir_weight[132][35],
reservoir_weight[132][36],
reservoir_weight[132][37],
reservoir_weight[132][38],
reservoir_weight[132][39],
reservoir_weight[132][40],
reservoir_weight[132][41],
reservoir_weight[132][42],
reservoir_weight[132][43],
reservoir_weight[132][44],
reservoir_weight[132][45],
reservoir_weight[132][46],
reservoir_weight[132][47],
reservoir_weight[132][48],
reservoir_weight[132][49],
reservoir_weight[132][50],
reservoir_weight[132][51],
reservoir_weight[132][52],
reservoir_weight[132][53],
reservoir_weight[132][54],
reservoir_weight[132][55],
reservoir_weight[132][56],
reservoir_weight[132][57],
reservoir_weight[132][58],
reservoir_weight[132][59],
reservoir_weight[132][60],
reservoir_weight[132][61],
reservoir_weight[132][62],
reservoir_weight[132][63],
reservoir_weight[132][64],
reservoir_weight[132][65],
reservoir_weight[132][66],
reservoir_weight[132][67],
reservoir_weight[132][68],
reservoir_weight[132][69],
reservoir_weight[132][70],
reservoir_weight[132][71],
reservoir_weight[132][72],
reservoir_weight[132][73],
reservoir_weight[132][74],
reservoir_weight[132][75],
reservoir_weight[132][76],
reservoir_weight[132][77],
reservoir_weight[132][78],
reservoir_weight[132][79],
reservoir_weight[132][80],
reservoir_weight[132][81],
reservoir_weight[132][82],
reservoir_weight[132][83],
reservoir_weight[132][84],
reservoir_weight[132][85],
reservoir_weight[132][86],
reservoir_weight[132][87],
reservoir_weight[132][88],
reservoir_weight[132][89],
reservoir_weight[132][90],
reservoir_weight[132][91],
reservoir_weight[132][92],
reservoir_weight[132][93],
reservoir_weight[132][94],
reservoir_weight[132][95],
reservoir_weight[132][96],
reservoir_weight[132][97],
reservoir_weight[132][98],
reservoir_weight[132][99],
reservoir_weight[132][100],
reservoir_weight[132][101],
reservoir_weight[132][102],
reservoir_weight[132][103],
reservoir_weight[132][104],
reservoir_weight[132][105],
reservoir_weight[132][106],
reservoir_weight[132][107],
reservoir_weight[132][108],
reservoir_weight[132][109],
reservoir_weight[132][110],
reservoir_weight[132][111],
reservoir_weight[132][112],
reservoir_weight[132][113],
reservoir_weight[132][114],
reservoir_weight[132][115],
reservoir_weight[132][116],
reservoir_weight[132][117],
reservoir_weight[132][118],
reservoir_weight[132][119],
reservoir_weight[132][120],
reservoir_weight[132][121],
reservoir_weight[132][122],
reservoir_weight[132][123],
reservoir_weight[132][124],
reservoir_weight[132][125],
reservoir_weight[132][126],
reservoir_weight[132][127],
reservoir_weight[132][128],
reservoir_weight[132][129],
reservoir_weight[132][130],
reservoir_weight[132][131],
reservoir_weight[132][132],
reservoir_weight[132][133],
reservoir_weight[132][134],
reservoir_weight[132][135],
reservoir_weight[132][136],
reservoir_weight[132][137],
reservoir_weight[132][138],
reservoir_weight[132][139],
reservoir_weight[132][140],
reservoir_weight[132][141],
reservoir_weight[132][142],
reservoir_weight[132][143],
reservoir_weight[132][144],
reservoir_weight[132][145],
reservoir_weight[132][146],
reservoir_weight[132][147],
reservoir_weight[132][148],
reservoir_weight[132][149],
reservoir_weight[132][150],
reservoir_weight[132][151],
reservoir_weight[132][152],
reservoir_weight[132][153],
reservoir_weight[132][154],
reservoir_weight[132][155],
reservoir_weight[132][156],
reservoir_weight[132][157],
reservoir_weight[132][158],
reservoir_weight[132][159],
reservoir_weight[132][160],
reservoir_weight[132][161],
reservoir_weight[132][162],
reservoir_weight[132][163],
reservoir_weight[132][164],
reservoir_weight[132][165],
reservoir_weight[132][166],
reservoir_weight[132][167],
reservoir_weight[132][168],
reservoir_weight[132][169],
reservoir_weight[132][170],
reservoir_weight[132][171],
reservoir_weight[132][172],
reservoir_weight[132][173],
reservoir_weight[132][174],
reservoir_weight[132][175],
reservoir_weight[132][176],
reservoir_weight[132][177],
reservoir_weight[132][178],
reservoir_weight[132][179],
reservoir_weight[132][180],
reservoir_weight[132][181],
reservoir_weight[132][182],
reservoir_weight[132][183],
reservoir_weight[132][184],
reservoir_weight[132][185],
reservoir_weight[132][186],
reservoir_weight[132][187],
reservoir_weight[132][188],
reservoir_weight[132][189],
reservoir_weight[132][190],
reservoir_weight[132][191],
reservoir_weight[132][192],
reservoir_weight[132][193],
reservoir_weight[132][194],
reservoir_weight[132][195],
reservoir_weight[132][196],
reservoir_weight[132][197],
reservoir_weight[132][198],
reservoir_weight[132][199]
},
{reservoir_weight[133][0],
reservoir_weight[133][1],
reservoir_weight[133][2],
reservoir_weight[133][3],
reservoir_weight[133][4],
reservoir_weight[133][5],
reservoir_weight[133][6],
reservoir_weight[133][7],
reservoir_weight[133][8],
reservoir_weight[133][9],
reservoir_weight[133][10],
reservoir_weight[133][11],
reservoir_weight[133][12],
reservoir_weight[133][13],
reservoir_weight[133][14],
reservoir_weight[133][15],
reservoir_weight[133][16],
reservoir_weight[133][17],
reservoir_weight[133][18],
reservoir_weight[133][19],
reservoir_weight[133][20],
reservoir_weight[133][21],
reservoir_weight[133][22],
reservoir_weight[133][23],
reservoir_weight[133][24],
reservoir_weight[133][25],
reservoir_weight[133][26],
reservoir_weight[133][27],
reservoir_weight[133][28],
reservoir_weight[133][29],
reservoir_weight[133][30],
reservoir_weight[133][31],
reservoir_weight[133][32],
reservoir_weight[133][33],
reservoir_weight[133][34],
reservoir_weight[133][35],
reservoir_weight[133][36],
reservoir_weight[133][37],
reservoir_weight[133][38],
reservoir_weight[133][39],
reservoir_weight[133][40],
reservoir_weight[133][41],
reservoir_weight[133][42],
reservoir_weight[133][43],
reservoir_weight[133][44],
reservoir_weight[133][45],
reservoir_weight[133][46],
reservoir_weight[133][47],
reservoir_weight[133][48],
reservoir_weight[133][49],
reservoir_weight[133][50],
reservoir_weight[133][51],
reservoir_weight[133][52],
reservoir_weight[133][53],
reservoir_weight[133][54],
reservoir_weight[133][55],
reservoir_weight[133][56],
reservoir_weight[133][57],
reservoir_weight[133][58],
reservoir_weight[133][59],
reservoir_weight[133][60],
reservoir_weight[133][61],
reservoir_weight[133][62],
reservoir_weight[133][63],
reservoir_weight[133][64],
reservoir_weight[133][65],
reservoir_weight[133][66],
reservoir_weight[133][67],
reservoir_weight[133][68],
reservoir_weight[133][69],
reservoir_weight[133][70],
reservoir_weight[133][71],
reservoir_weight[133][72],
reservoir_weight[133][73],
reservoir_weight[133][74],
reservoir_weight[133][75],
reservoir_weight[133][76],
reservoir_weight[133][77],
reservoir_weight[133][78],
reservoir_weight[133][79],
reservoir_weight[133][80],
reservoir_weight[133][81],
reservoir_weight[133][82],
reservoir_weight[133][83],
reservoir_weight[133][84],
reservoir_weight[133][85],
reservoir_weight[133][86],
reservoir_weight[133][87],
reservoir_weight[133][88],
reservoir_weight[133][89],
reservoir_weight[133][90],
reservoir_weight[133][91],
reservoir_weight[133][92],
reservoir_weight[133][93],
reservoir_weight[133][94],
reservoir_weight[133][95],
reservoir_weight[133][96],
reservoir_weight[133][97],
reservoir_weight[133][98],
reservoir_weight[133][99],
reservoir_weight[133][100],
reservoir_weight[133][101],
reservoir_weight[133][102],
reservoir_weight[133][103],
reservoir_weight[133][104],
reservoir_weight[133][105],
reservoir_weight[133][106],
reservoir_weight[133][107],
reservoir_weight[133][108],
reservoir_weight[133][109],
reservoir_weight[133][110],
reservoir_weight[133][111],
reservoir_weight[133][112],
reservoir_weight[133][113],
reservoir_weight[133][114],
reservoir_weight[133][115],
reservoir_weight[133][116],
reservoir_weight[133][117],
reservoir_weight[133][118],
reservoir_weight[133][119],
reservoir_weight[133][120],
reservoir_weight[133][121],
reservoir_weight[133][122],
reservoir_weight[133][123],
reservoir_weight[133][124],
reservoir_weight[133][125],
reservoir_weight[133][126],
reservoir_weight[133][127],
reservoir_weight[133][128],
reservoir_weight[133][129],
reservoir_weight[133][130],
reservoir_weight[133][131],
reservoir_weight[133][132],
reservoir_weight[133][133],
reservoir_weight[133][134],
reservoir_weight[133][135],
reservoir_weight[133][136],
reservoir_weight[133][137],
reservoir_weight[133][138],
reservoir_weight[133][139],
reservoir_weight[133][140],
reservoir_weight[133][141],
reservoir_weight[133][142],
reservoir_weight[133][143],
reservoir_weight[133][144],
reservoir_weight[133][145],
reservoir_weight[133][146],
reservoir_weight[133][147],
reservoir_weight[133][148],
reservoir_weight[133][149],
reservoir_weight[133][150],
reservoir_weight[133][151],
reservoir_weight[133][152],
reservoir_weight[133][153],
reservoir_weight[133][154],
reservoir_weight[133][155],
reservoir_weight[133][156],
reservoir_weight[133][157],
reservoir_weight[133][158],
reservoir_weight[133][159],
reservoir_weight[133][160],
reservoir_weight[133][161],
reservoir_weight[133][162],
reservoir_weight[133][163],
reservoir_weight[133][164],
reservoir_weight[133][165],
reservoir_weight[133][166],
reservoir_weight[133][167],
reservoir_weight[133][168],
reservoir_weight[133][169],
reservoir_weight[133][170],
reservoir_weight[133][171],
reservoir_weight[133][172],
reservoir_weight[133][173],
reservoir_weight[133][174],
reservoir_weight[133][175],
reservoir_weight[133][176],
reservoir_weight[133][177],
reservoir_weight[133][178],
reservoir_weight[133][179],
reservoir_weight[133][180],
reservoir_weight[133][181],
reservoir_weight[133][182],
reservoir_weight[133][183],
reservoir_weight[133][184],
reservoir_weight[133][185],
reservoir_weight[133][186],
reservoir_weight[133][187],
reservoir_weight[133][188],
reservoir_weight[133][189],
reservoir_weight[133][190],
reservoir_weight[133][191],
reservoir_weight[133][192],
reservoir_weight[133][193],
reservoir_weight[133][194],
reservoir_weight[133][195],
reservoir_weight[133][196],
reservoir_weight[133][197],
reservoir_weight[133][198],
reservoir_weight[133][199]
},
{reservoir_weight[134][0],
reservoir_weight[134][1],
reservoir_weight[134][2],
reservoir_weight[134][3],
reservoir_weight[134][4],
reservoir_weight[134][5],
reservoir_weight[134][6],
reservoir_weight[134][7],
reservoir_weight[134][8],
reservoir_weight[134][9],
reservoir_weight[134][10],
reservoir_weight[134][11],
reservoir_weight[134][12],
reservoir_weight[134][13],
reservoir_weight[134][14],
reservoir_weight[134][15],
reservoir_weight[134][16],
reservoir_weight[134][17],
reservoir_weight[134][18],
reservoir_weight[134][19],
reservoir_weight[134][20],
reservoir_weight[134][21],
reservoir_weight[134][22],
reservoir_weight[134][23],
reservoir_weight[134][24],
reservoir_weight[134][25],
reservoir_weight[134][26],
reservoir_weight[134][27],
reservoir_weight[134][28],
reservoir_weight[134][29],
reservoir_weight[134][30],
reservoir_weight[134][31],
reservoir_weight[134][32],
reservoir_weight[134][33],
reservoir_weight[134][34],
reservoir_weight[134][35],
reservoir_weight[134][36],
reservoir_weight[134][37],
reservoir_weight[134][38],
reservoir_weight[134][39],
reservoir_weight[134][40],
reservoir_weight[134][41],
reservoir_weight[134][42],
reservoir_weight[134][43],
reservoir_weight[134][44],
reservoir_weight[134][45],
reservoir_weight[134][46],
reservoir_weight[134][47],
reservoir_weight[134][48],
reservoir_weight[134][49],
reservoir_weight[134][50],
reservoir_weight[134][51],
reservoir_weight[134][52],
reservoir_weight[134][53],
reservoir_weight[134][54],
reservoir_weight[134][55],
reservoir_weight[134][56],
reservoir_weight[134][57],
reservoir_weight[134][58],
reservoir_weight[134][59],
reservoir_weight[134][60],
reservoir_weight[134][61],
reservoir_weight[134][62],
reservoir_weight[134][63],
reservoir_weight[134][64],
reservoir_weight[134][65],
reservoir_weight[134][66],
reservoir_weight[134][67],
reservoir_weight[134][68],
reservoir_weight[134][69],
reservoir_weight[134][70],
reservoir_weight[134][71],
reservoir_weight[134][72],
reservoir_weight[134][73],
reservoir_weight[134][74],
reservoir_weight[134][75],
reservoir_weight[134][76],
reservoir_weight[134][77],
reservoir_weight[134][78],
reservoir_weight[134][79],
reservoir_weight[134][80],
reservoir_weight[134][81],
reservoir_weight[134][82],
reservoir_weight[134][83],
reservoir_weight[134][84],
reservoir_weight[134][85],
reservoir_weight[134][86],
reservoir_weight[134][87],
reservoir_weight[134][88],
reservoir_weight[134][89],
reservoir_weight[134][90],
reservoir_weight[134][91],
reservoir_weight[134][92],
reservoir_weight[134][93],
reservoir_weight[134][94],
reservoir_weight[134][95],
reservoir_weight[134][96],
reservoir_weight[134][97],
reservoir_weight[134][98],
reservoir_weight[134][99],
reservoir_weight[134][100],
reservoir_weight[134][101],
reservoir_weight[134][102],
reservoir_weight[134][103],
reservoir_weight[134][104],
reservoir_weight[134][105],
reservoir_weight[134][106],
reservoir_weight[134][107],
reservoir_weight[134][108],
reservoir_weight[134][109],
reservoir_weight[134][110],
reservoir_weight[134][111],
reservoir_weight[134][112],
reservoir_weight[134][113],
reservoir_weight[134][114],
reservoir_weight[134][115],
reservoir_weight[134][116],
reservoir_weight[134][117],
reservoir_weight[134][118],
reservoir_weight[134][119],
reservoir_weight[134][120],
reservoir_weight[134][121],
reservoir_weight[134][122],
reservoir_weight[134][123],
reservoir_weight[134][124],
reservoir_weight[134][125],
reservoir_weight[134][126],
reservoir_weight[134][127],
reservoir_weight[134][128],
reservoir_weight[134][129],
reservoir_weight[134][130],
reservoir_weight[134][131],
reservoir_weight[134][132],
reservoir_weight[134][133],
reservoir_weight[134][134],
reservoir_weight[134][135],
reservoir_weight[134][136],
reservoir_weight[134][137],
reservoir_weight[134][138],
reservoir_weight[134][139],
reservoir_weight[134][140],
reservoir_weight[134][141],
reservoir_weight[134][142],
reservoir_weight[134][143],
reservoir_weight[134][144],
reservoir_weight[134][145],
reservoir_weight[134][146],
reservoir_weight[134][147],
reservoir_weight[134][148],
reservoir_weight[134][149],
reservoir_weight[134][150],
reservoir_weight[134][151],
reservoir_weight[134][152],
reservoir_weight[134][153],
reservoir_weight[134][154],
reservoir_weight[134][155],
reservoir_weight[134][156],
reservoir_weight[134][157],
reservoir_weight[134][158],
reservoir_weight[134][159],
reservoir_weight[134][160],
reservoir_weight[134][161],
reservoir_weight[134][162],
reservoir_weight[134][163],
reservoir_weight[134][164],
reservoir_weight[134][165],
reservoir_weight[134][166],
reservoir_weight[134][167],
reservoir_weight[134][168],
reservoir_weight[134][169],
reservoir_weight[134][170],
reservoir_weight[134][171],
reservoir_weight[134][172],
reservoir_weight[134][173],
reservoir_weight[134][174],
reservoir_weight[134][175],
reservoir_weight[134][176],
reservoir_weight[134][177],
reservoir_weight[134][178],
reservoir_weight[134][179],
reservoir_weight[134][180],
reservoir_weight[134][181],
reservoir_weight[134][182],
reservoir_weight[134][183],
reservoir_weight[134][184],
reservoir_weight[134][185],
reservoir_weight[134][186],
reservoir_weight[134][187],
reservoir_weight[134][188],
reservoir_weight[134][189],
reservoir_weight[134][190],
reservoir_weight[134][191],
reservoir_weight[134][192],
reservoir_weight[134][193],
reservoir_weight[134][194],
reservoir_weight[134][195],
reservoir_weight[134][196],
reservoir_weight[134][197],
reservoir_weight[134][198],
reservoir_weight[134][199]
},
{reservoir_weight[135][0],
reservoir_weight[135][1],
reservoir_weight[135][2],
reservoir_weight[135][3],
reservoir_weight[135][4],
reservoir_weight[135][5],
reservoir_weight[135][6],
reservoir_weight[135][7],
reservoir_weight[135][8],
reservoir_weight[135][9],
reservoir_weight[135][10],
reservoir_weight[135][11],
reservoir_weight[135][12],
reservoir_weight[135][13],
reservoir_weight[135][14],
reservoir_weight[135][15],
reservoir_weight[135][16],
reservoir_weight[135][17],
reservoir_weight[135][18],
reservoir_weight[135][19],
reservoir_weight[135][20],
reservoir_weight[135][21],
reservoir_weight[135][22],
reservoir_weight[135][23],
reservoir_weight[135][24],
reservoir_weight[135][25],
reservoir_weight[135][26],
reservoir_weight[135][27],
reservoir_weight[135][28],
reservoir_weight[135][29],
reservoir_weight[135][30],
reservoir_weight[135][31],
reservoir_weight[135][32],
reservoir_weight[135][33],
reservoir_weight[135][34],
reservoir_weight[135][35],
reservoir_weight[135][36],
reservoir_weight[135][37],
reservoir_weight[135][38],
reservoir_weight[135][39],
reservoir_weight[135][40],
reservoir_weight[135][41],
reservoir_weight[135][42],
reservoir_weight[135][43],
reservoir_weight[135][44],
reservoir_weight[135][45],
reservoir_weight[135][46],
reservoir_weight[135][47],
reservoir_weight[135][48],
reservoir_weight[135][49],
reservoir_weight[135][50],
reservoir_weight[135][51],
reservoir_weight[135][52],
reservoir_weight[135][53],
reservoir_weight[135][54],
reservoir_weight[135][55],
reservoir_weight[135][56],
reservoir_weight[135][57],
reservoir_weight[135][58],
reservoir_weight[135][59],
reservoir_weight[135][60],
reservoir_weight[135][61],
reservoir_weight[135][62],
reservoir_weight[135][63],
reservoir_weight[135][64],
reservoir_weight[135][65],
reservoir_weight[135][66],
reservoir_weight[135][67],
reservoir_weight[135][68],
reservoir_weight[135][69],
reservoir_weight[135][70],
reservoir_weight[135][71],
reservoir_weight[135][72],
reservoir_weight[135][73],
reservoir_weight[135][74],
reservoir_weight[135][75],
reservoir_weight[135][76],
reservoir_weight[135][77],
reservoir_weight[135][78],
reservoir_weight[135][79],
reservoir_weight[135][80],
reservoir_weight[135][81],
reservoir_weight[135][82],
reservoir_weight[135][83],
reservoir_weight[135][84],
reservoir_weight[135][85],
reservoir_weight[135][86],
reservoir_weight[135][87],
reservoir_weight[135][88],
reservoir_weight[135][89],
reservoir_weight[135][90],
reservoir_weight[135][91],
reservoir_weight[135][92],
reservoir_weight[135][93],
reservoir_weight[135][94],
reservoir_weight[135][95],
reservoir_weight[135][96],
reservoir_weight[135][97],
reservoir_weight[135][98],
reservoir_weight[135][99],
reservoir_weight[135][100],
reservoir_weight[135][101],
reservoir_weight[135][102],
reservoir_weight[135][103],
reservoir_weight[135][104],
reservoir_weight[135][105],
reservoir_weight[135][106],
reservoir_weight[135][107],
reservoir_weight[135][108],
reservoir_weight[135][109],
reservoir_weight[135][110],
reservoir_weight[135][111],
reservoir_weight[135][112],
reservoir_weight[135][113],
reservoir_weight[135][114],
reservoir_weight[135][115],
reservoir_weight[135][116],
reservoir_weight[135][117],
reservoir_weight[135][118],
reservoir_weight[135][119],
reservoir_weight[135][120],
reservoir_weight[135][121],
reservoir_weight[135][122],
reservoir_weight[135][123],
reservoir_weight[135][124],
reservoir_weight[135][125],
reservoir_weight[135][126],
reservoir_weight[135][127],
reservoir_weight[135][128],
reservoir_weight[135][129],
reservoir_weight[135][130],
reservoir_weight[135][131],
reservoir_weight[135][132],
reservoir_weight[135][133],
reservoir_weight[135][134],
reservoir_weight[135][135],
reservoir_weight[135][136],
reservoir_weight[135][137],
reservoir_weight[135][138],
reservoir_weight[135][139],
reservoir_weight[135][140],
reservoir_weight[135][141],
reservoir_weight[135][142],
reservoir_weight[135][143],
reservoir_weight[135][144],
reservoir_weight[135][145],
reservoir_weight[135][146],
reservoir_weight[135][147],
reservoir_weight[135][148],
reservoir_weight[135][149],
reservoir_weight[135][150],
reservoir_weight[135][151],
reservoir_weight[135][152],
reservoir_weight[135][153],
reservoir_weight[135][154],
reservoir_weight[135][155],
reservoir_weight[135][156],
reservoir_weight[135][157],
reservoir_weight[135][158],
reservoir_weight[135][159],
reservoir_weight[135][160],
reservoir_weight[135][161],
reservoir_weight[135][162],
reservoir_weight[135][163],
reservoir_weight[135][164],
reservoir_weight[135][165],
reservoir_weight[135][166],
reservoir_weight[135][167],
reservoir_weight[135][168],
reservoir_weight[135][169],
reservoir_weight[135][170],
reservoir_weight[135][171],
reservoir_weight[135][172],
reservoir_weight[135][173],
reservoir_weight[135][174],
reservoir_weight[135][175],
reservoir_weight[135][176],
reservoir_weight[135][177],
reservoir_weight[135][178],
reservoir_weight[135][179],
reservoir_weight[135][180],
reservoir_weight[135][181],
reservoir_weight[135][182],
reservoir_weight[135][183],
reservoir_weight[135][184],
reservoir_weight[135][185],
reservoir_weight[135][186],
reservoir_weight[135][187],
reservoir_weight[135][188],
reservoir_weight[135][189],
reservoir_weight[135][190],
reservoir_weight[135][191],
reservoir_weight[135][192],
reservoir_weight[135][193],
reservoir_weight[135][194],
reservoir_weight[135][195],
reservoir_weight[135][196],
reservoir_weight[135][197],
reservoir_weight[135][198],
reservoir_weight[135][199]
},
{reservoir_weight[136][0],
reservoir_weight[136][1],
reservoir_weight[136][2],
reservoir_weight[136][3],
reservoir_weight[136][4],
reservoir_weight[136][5],
reservoir_weight[136][6],
reservoir_weight[136][7],
reservoir_weight[136][8],
reservoir_weight[136][9],
reservoir_weight[136][10],
reservoir_weight[136][11],
reservoir_weight[136][12],
reservoir_weight[136][13],
reservoir_weight[136][14],
reservoir_weight[136][15],
reservoir_weight[136][16],
reservoir_weight[136][17],
reservoir_weight[136][18],
reservoir_weight[136][19],
reservoir_weight[136][20],
reservoir_weight[136][21],
reservoir_weight[136][22],
reservoir_weight[136][23],
reservoir_weight[136][24],
reservoir_weight[136][25],
reservoir_weight[136][26],
reservoir_weight[136][27],
reservoir_weight[136][28],
reservoir_weight[136][29],
reservoir_weight[136][30],
reservoir_weight[136][31],
reservoir_weight[136][32],
reservoir_weight[136][33],
reservoir_weight[136][34],
reservoir_weight[136][35],
reservoir_weight[136][36],
reservoir_weight[136][37],
reservoir_weight[136][38],
reservoir_weight[136][39],
reservoir_weight[136][40],
reservoir_weight[136][41],
reservoir_weight[136][42],
reservoir_weight[136][43],
reservoir_weight[136][44],
reservoir_weight[136][45],
reservoir_weight[136][46],
reservoir_weight[136][47],
reservoir_weight[136][48],
reservoir_weight[136][49],
reservoir_weight[136][50],
reservoir_weight[136][51],
reservoir_weight[136][52],
reservoir_weight[136][53],
reservoir_weight[136][54],
reservoir_weight[136][55],
reservoir_weight[136][56],
reservoir_weight[136][57],
reservoir_weight[136][58],
reservoir_weight[136][59],
reservoir_weight[136][60],
reservoir_weight[136][61],
reservoir_weight[136][62],
reservoir_weight[136][63],
reservoir_weight[136][64],
reservoir_weight[136][65],
reservoir_weight[136][66],
reservoir_weight[136][67],
reservoir_weight[136][68],
reservoir_weight[136][69],
reservoir_weight[136][70],
reservoir_weight[136][71],
reservoir_weight[136][72],
reservoir_weight[136][73],
reservoir_weight[136][74],
reservoir_weight[136][75],
reservoir_weight[136][76],
reservoir_weight[136][77],
reservoir_weight[136][78],
reservoir_weight[136][79],
reservoir_weight[136][80],
reservoir_weight[136][81],
reservoir_weight[136][82],
reservoir_weight[136][83],
reservoir_weight[136][84],
reservoir_weight[136][85],
reservoir_weight[136][86],
reservoir_weight[136][87],
reservoir_weight[136][88],
reservoir_weight[136][89],
reservoir_weight[136][90],
reservoir_weight[136][91],
reservoir_weight[136][92],
reservoir_weight[136][93],
reservoir_weight[136][94],
reservoir_weight[136][95],
reservoir_weight[136][96],
reservoir_weight[136][97],
reservoir_weight[136][98],
reservoir_weight[136][99],
reservoir_weight[136][100],
reservoir_weight[136][101],
reservoir_weight[136][102],
reservoir_weight[136][103],
reservoir_weight[136][104],
reservoir_weight[136][105],
reservoir_weight[136][106],
reservoir_weight[136][107],
reservoir_weight[136][108],
reservoir_weight[136][109],
reservoir_weight[136][110],
reservoir_weight[136][111],
reservoir_weight[136][112],
reservoir_weight[136][113],
reservoir_weight[136][114],
reservoir_weight[136][115],
reservoir_weight[136][116],
reservoir_weight[136][117],
reservoir_weight[136][118],
reservoir_weight[136][119],
reservoir_weight[136][120],
reservoir_weight[136][121],
reservoir_weight[136][122],
reservoir_weight[136][123],
reservoir_weight[136][124],
reservoir_weight[136][125],
reservoir_weight[136][126],
reservoir_weight[136][127],
reservoir_weight[136][128],
reservoir_weight[136][129],
reservoir_weight[136][130],
reservoir_weight[136][131],
reservoir_weight[136][132],
reservoir_weight[136][133],
reservoir_weight[136][134],
reservoir_weight[136][135],
reservoir_weight[136][136],
reservoir_weight[136][137],
reservoir_weight[136][138],
reservoir_weight[136][139],
reservoir_weight[136][140],
reservoir_weight[136][141],
reservoir_weight[136][142],
reservoir_weight[136][143],
reservoir_weight[136][144],
reservoir_weight[136][145],
reservoir_weight[136][146],
reservoir_weight[136][147],
reservoir_weight[136][148],
reservoir_weight[136][149],
reservoir_weight[136][150],
reservoir_weight[136][151],
reservoir_weight[136][152],
reservoir_weight[136][153],
reservoir_weight[136][154],
reservoir_weight[136][155],
reservoir_weight[136][156],
reservoir_weight[136][157],
reservoir_weight[136][158],
reservoir_weight[136][159],
reservoir_weight[136][160],
reservoir_weight[136][161],
reservoir_weight[136][162],
reservoir_weight[136][163],
reservoir_weight[136][164],
reservoir_weight[136][165],
reservoir_weight[136][166],
reservoir_weight[136][167],
reservoir_weight[136][168],
reservoir_weight[136][169],
reservoir_weight[136][170],
reservoir_weight[136][171],
reservoir_weight[136][172],
reservoir_weight[136][173],
reservoir_weight[136][174],
reservoir_weight[136][175],
reservoir_weight[136][176],
reservoir_weight[136][177],
reservoir_weight[136][178],
reservoir_weight[136][179],
reservoir_weight[136][180],
reservoir_weight[136][181],
reservoir_weight[136][182],
reservoir_weight[136][183],
reservoir_weight[136][184],
reservoir_weight[136][185],
reservoir_weight[136][186],
reservoir_weight[136][187],
reservoir_weight[136][188],
reservoir_weight[136][189],
reservoir_weight[136][190],
reservoir_weight[136][191],
reservoir_weight[136][192],
reservoir_weight[136][193],
reservoir_weight[136][194],
reservoir_weight[136][195],
reservoir_weight[136][196],
reservoir_weight[136][197],
reservoir_weight[136][198],
reservoir_weight[136][199]
},
{reservoir_weight[137][0],
reservoir_weight[137][1],
reservoir_weight[137][2],
reservoir_weight[137][3],
reservoir_weight[137][4],
reservoir_weight[137][5],
reservoir_weight[137][6],
reservoir_weight[137][7],
reservoir_weight[137][8],
reservoir_weight[137][9],
reservoir_weight[137][10],
reservoir_weight[137][11],
reservoir_weight[137][12],
reservoir_weight[137][13],
reservoir_weight[137][14],
reservoir_weight[137][15],
reservoir_weight[137][16],
reservoir_weight[137][17],
reservoir_weight[137][18],
reservoir_weight[137][19],
reservoir_weight[137][20],
reservoir_weight[137][21],
reservoir_weight[137][22],
reservoir_weight[137][23],
reservoir_weight[137][24],
reservoir_weight[137][25],
reservoir_weight[137][26],
reservoir_weight[137][27],
reservoir_weight[137][28],
reservoir_weight[137][29],
reservoir_weight[137][30],
reservoir_weight[137][31],
reservoir_weight[137][32],
reservoir_weight[137][33],
reservoir_weight[137][34],
reservoir_weight[137][35],
reservoir_weight[137][36],
reservoir_weight[137][37],
reservoir_weight[137][38],
reservoir_weight[137][39],
reservoir_weight[137][40],
reservoir_weight[137][41],
reservoir_weight[137][42],
reservoir_weight[137][43],
reservoir_weight[137][44],
reservoir_weight[137][45],
reservoir_weight[137][46],
reservoir_weight[137][47],
reservoir_weight[137][48],
reservoir_weight[137][49],
reservoir_weight[137][50],
reservoir_weight[137][51],
reservoir_weight[137][52],
reservoir_weight[137][53],
reservoir_weight[137][54],
reservoir_weight[137][55],
reservoir_weight[137][56],
reservoir_weight[137][57],
reservoir_weight[137][58],
reservoir_weight[137][59],
reservoir_weight[137][60],
reservoir_weight[137][61],
reservoir_weight[137][62],
reservoir_weight[137][63],
reservoir_weight[137][64],
reservoir_weight[137][65],
reservoir_weight[137][66],
reservoir_weight[137][67],
reservoir_weight[137][68],
reservoir_weight[137][69],
reservoir_weight[137][70],
reservoir_weight[137][71],
reservoir_weight[137][72],
reservoir_weight[137][73],
reservoir_weight[137][74],
reservoir_weight[137][75],
reservoir_weight[137][76],
reservoir_weight[137][77],
reservoir_weight[137][78],
reservoir_weight[137][79],
reservoir_weight[137][80],
reservoir_weight[137][81],
reservoir_weight[137][82],
reservoir_weight[137][83],
reservoir_weight[137][84],
reservoir_weight[137][85],
reservoir_weight[137][86],
reservoir_weight[137][87],
reservoir_weight[137][88],
reservoir_weight[137][89],
reservoir_weight[137][90],
reservoir_weight[137][91],
reservoir_weight[137][92],
reservoir_weight[137][93],
reservoir_weight[137][94],
reservoir_weight[137][95],
reservoir_weight[137][96],
reservoir_weight[137][97],
reservoir_weight[137][98],
reservoir_weight[137][99],
reservoir_weight[137][100],
reservoir_weight[137][101],
reservoir_weight[137][102],
reservoir_weight[137][103],
reservoir_weight[137][104],
reservoir_weight[137][105],
reservoir_weight[137][106],
reservoir_weight[137][107],
reservoir_weight[137][108],
reservoir_weight[137][109],
reservoir_weight[137][110],
reservoir_weight[137][111],
reservoir_weight[137][112],
reservoir_weight[137][113],
reservoir_weight[137][114],
reservoir_weight[137][115],
reservoir_weight[137][116],
reservoir_weight[137][117],
reservoir_weight[137][118],
reservoir_weight[137][119],
reservoir_weight[137][120],
reservoir_weight[137][121],
reservoir_weight[137][122],
reservoir_weight[137][123],
reservoir_weight[137][124],
reservoir_weight[137][125],
reservoir_weight[137][126],
reservoir_weight[137][127],
reservoir_weight[137][128],
reservoir_weight[137][129],
reservoir_weight[137][130],
reservoir_weight[137][131],
reservoir_weight[137][132],
reservoir_weight[137][133],
reservoir_weight[137][134],
reservoir_weight[137][135],
reservoir_weight[137][136],
reservoir_weight[137][137],
reservoir_weight[137][138],
reservoir_weight[137][139],
reservoir_weight[137][140],
reservoir_weight[137][141],
reservoir_weight[137][142],
reservoir_weight[137][143],
reservoir_weight[137][144],
reservoir_weight[137][145],
reservoir_weight[137][146],
reservoir_weight[137][147],
reservoir_weight[137][148],
reservoir_weight[137][149],
reservoir_weight[137][150],
reservoir_weight[137][151],
reservoir_weight[137][152],
reservoir_weight[137][153],
reservoir_weight[137][154],
reservoir_weight[137][155],
reservoir_weight[137][156],
reservoir_weight[137][157],
reservoir_weight[137][158],
reservoir_weight[137][159],
reservoir_weight[137][160],
reservoir_weight[137][161],
reservoir_weight[137][162],
reservoir_weight[137][163],
reservoir_weight[137][164],
reservoir_weight[137][165],
reservoir_weight[137][166],
reservoir_weight[137][167],
reservoir_weight[137][168],
reservoir_weight[137][169],
reservoir_weight[137][170],
reservoir_weight[137][171],
reservoir_weight[137][172],
reservoir_weight[137][173],
reservoir_weight[137][174],
reservoir_weight[137][175],
reservoir_weight[137][176],
reservoir_weight[137][177],
reservoir_weight[137][178],
reservoir_weight[137][179],
reservoir_weight[137][180],
reservoir_weight[137][181],
reservoir_weight[137][182],
reservoir_weight[137][183],
reservoir_weight[137][184],
reservoir_weight[137][185],
reservoir_weight[137][186],
reservoir_weight[137][187],
reservoir_weight[137][188],
reservoir_weight[137][189],
reservoir_weight[137][190],
reservoir_weight[137][191],
reservoir_weight[137][192],
reservoir_weight[137][193],
reservoir_weight[137][194],
reservoir_weight[137][195],
reservoir_weight[137][196],
reservoir_weight[137][197],
reservoir_weight[137][198],
reservoir_weight[137][199]
},
{reservoir_weight[138][0],
reservoir_weight[138][1],
reservoir_weight[138][2],
reservoir_weight[138][3],
reservoir_weight[138][4],
reservoir_weight[138][5],
reservoir_weight[138][6],
reservoir_weight[138][7],
reservoir_weight[138][8],
reservoir_weight[138][9],
reservoir_weight[138][10],
reservoir_weight[138][11],
reservoir_weight[138][12],
reservoir_weight[138][13],
reservoir_weight[138][14],
reservoir_weight[138][15],
reservoir_weight[138][16],
reservoir_weight[138][17],
reservoir_weight[138][18],
reservoir_weight[138][19],
reservoir_weight[138][20],
reservoir_weight[138][21],
reservoir_weight[138][22],
reservoir_weight[138][23],
reservoir_weight[138][24],
reservoir_weight[138][25],
reservoir_weight[138][26],
reservoir_weight[138][27],
reservoir_weight[138][28],
reservoir_weight[138][29],
reservoir_weight[138][30],
reservoir_weight[138][31],
reservoir_weight[138][32],
reservoir_weight[138][33],
reservoir_weight[138][34],
reservoir_weight[138][35],
reservoir_weight[138][36],
reservoir_weight[138][37],
reservoir_weight[138][38],
reservoir_weight[138][39],
reservoir_weight[138][40],
reservoir_weight[138][41],
reservoir_weight[138][42],
reservoir_weight[138][43],
reservoir_weight[138][44],
reservoir_weight[138][45],
reservoir_weight[138][46],
reservoir_weight[138][47],
reservoir_weight[138][48],
reservoir_weight[138][49],
reservoir_weight[138][50],
reservoir_weight[138][51],
reservoir_weight[138][52],
reservoir_weight[138][53],
reservoir_weight[138][54],
reservoir_weight[138][55],
reservoir_weight[138][56],
reservoir_weight[138][57],
reservoir_weight[138][58],
reservoir_weight[138][59],
reservoir_weight[138][60],
reservoir_weight[138][61],
reservoir_weight[138][62],
reservoir_weight[138][63],
reservoir_weight[138][64],
reservoir_weight[138][65],
reservoir_weight[138][66],
reservoir_weight[138][67],
reservoir_weight[138][68],
reservoir_weight[138][69],
reservoir_weight[138][70],
reservoir_weight[138][71],
reservoir_weight[138][72],
reservoir_weight[138][73],
reservoir_weight[138][74],
reservoir_weight[138][75],
reservoir_weight[138][76],
reservoir_weight[138][77],
reservoir_weight[138][78],
reservoir_weight[138][79],
reservoir_weight[138][80],
reservoir_weight[138][81],
reservoir_weight[138][82],
reservoir_weight[138][83],
reservoir_weight[138][84],
reservoir_weight[138][85],
reservoir_weight[138][86],
reservoir_weight[138][87],
reservoir_weight[138][88],
reservoir_weight[138][89],
reservoir_weight[138][90],
reservoir_weight[138][91],
reservoir_weight[138][92],
reservoir_weight[138][93],
reservoir_weight[138][94],
reservoir_weight[138][95],
reservoir_weight[138][96],
reservoir_weight[138][97],
reservoir_weight[138][98],
reservoir_weight[138][99],
reservoir_weight[138][100],
reservoir_weight[138][101],
reservoir_weight[138][102],
reservoir_weight[138][103],
reservoir_weight[138][104],
reservoir_weight[138][105],
reservoir_weight[138][106],
reservoir_weight[138][107],
reservoir_weight[138][108],
reservoir_weight[138][109],
reservoir_weight[138][110],
reservoir_weight[138][111],
reservoir_weight[138][112],
reservoir_weight[138][113],
reservoir_weight[138][114],
reservoir_weight[138][115],
reservoir_weight[138][116],
reservoir_weight[138][117],
reservoir_weight[138][118],
reservoir_weight[138][119],
reservoir_weight[138][120],
reservoir_weight[138][121],
reservoir_weight[138][122],
reservoir_weight[138][123],
reservoir_weight[138][124],
reservoir_weight[138][125],
reservoir_weight[138][126],
reservoir_weight[138][127],
reservoir_weight[138][128],
reservoir_weight[138][129],
reservoir_weight[138][130],
reservoir_weight[138][131],
reservoir_weight[138][132],
reservoir_weight[138][133],
reservoir_weight[138][134],
reservoir_weight[138][135],
reservoir_weight[138][136],
reservoir_weight[138][137],
reservoir_weight[138][138],
reservoir_weight[138][139],
reservoir_weight[138][140],
reservoir_weight[138][141],
reservoir_weight[138][142],
reservoir_weight[138][143],
reservoir_weight[138][144],
reservoir_weight[138][145],
reservoir_weight[138][146],
reservoir_weight[138][147],
reservoir_weight[138][148],
reservoir_weight[138][149],
reservoir_weight[138][150],
reservoir_weight[138][151],
reservoir_weight[138][152],
reservoir_weight[138][153],
reservoir_weight[138][154],
reservoir_weight[138][155],
reservoir_weight[138][156],
reservoir_weight[138][157],
reservoir_weight[138][158],
reservoir_weight[138][159],
reservoir_weight[138][160],
reservoir_weight[138][161],
reservoir_weight[138][162],
reservoir_weight[138][163],
reservoir_weight[138][164],
reservoir_weight[138][165],
reservoir_weight[138][166],
reservoir_weight[138][167],
reservoir_weight[138][168],
reservoir_weight[138][169],
reservoir_weight[138][170],
reservoir_weight[138][171],
reservoir_weight[138][172],
reservoir_weight[138][173],
reservoir_weight[138][174],
reservoir_weight[138][175],
reservoir_weight[138][176],
reservoir_weight[138][177],
reservoir_weight[138][178],
reservoir_weight[138][179],
reservoir_weight[138][180],
reservoir_weight[138][181],
reservoir_weight[138][182],
reservoir_weight[138][183],
reservoir_weight[138][184],
reservoir_weight[138][185],
reservoir_weight[138][186],
reservoir_weight[138][187],
reservoir_weight[138][188],
reservoir_weight[138][189],
reservoir_weight[138][190],
reservoir_weight[138][191],
reservoir_weight[138][192],
reservoir_weight[138][193],
reservoir_weight[138][194],
reservoir_weight[138][195],
reservoir_weight[138][196],
reservoir_weight[138][197],
reservoir_weight[138][198],
reservoir_weight[138][199]
},
{reservoir_weight[139][0],
reservoir_weight[139][1],
reservoir_weight[139][2],
reservoir_weight[139][3],
reservoir_weight[139][4],
reservoir_weight[139][5],
reservoir_weight[139][6],
reservoir_weight[139][7],
reservoir_weight[139][8],
reservoir_weight[139][9],
reservoir_weight[139][10],
reservoir_weight[139][11],
reservoir_weight[139][12],
reservoir_weight[139][13],
reservoir_weight[139][14],
reservoir_weight[139][15],
reservoir_weight[139][16],
reservoir_weight[139][17],
reservoir_weight[139][18],
reservoir_weight[139][19],
reservoir_weight[139][20],
reservoir_weight[139][21],
reservoir_weight[139][22],
reservoir_weight[139][23],
reservoir_weight[139][24],
reservoir_weight[139][25],
reservoir_weight[139][26],
reservoir_weight[139][27],
reservoir_weight[139][28],
reservoir_weight[139][29],
reservoir_weight[139][30],
reservoir_weight[139][31],
reservoir_weight[139][32],
reservoir_weight[139][33],
reservoir_weight[139][34],
reservoir_weight[139][35],
reservoir_weight[139][36],
reservoir_weight[139][37],
reservoir_weight[139][38],
reservoir_weight[139][39],
reservoir_weight[139][40],
reservoir_weight[139][41],
reservoir_weight[139][42],
reservoir_weight[139][43],
reservoir_weight[139][44],
reservoir_weight[139][45],
reservoir_weight[139][46],
reservoir_weight[139][47],
reservoir_weight[139][48],
reservoir_weight[139][49],
reservoir_weight[139][50],
reservoir_weight[139][51],
reservoir_weight[139][52],
reservoir_weight[139][53],
reservoir_weight[139][54],
reservoir_weight[139][55],
reservoir_weight[139][56],
reservoir_weight[139][57],
reservoir_weight[139][58],
reservoir_weight[139][59],
reservoir_weight[139][60],
reservoir_weight[139][61],
reservoir_weight[139][62],
reservoir_weight[139][63],
reservoir_weight[139][64],
reservoir_weight[139][65],
reservoir_weight[139][66],
reservoir_weight[139][67],
reservoir_weight[139][68],
reservoir_weight[139][69],
reservoir_weight[139][70],
reservoir_weight[139][71],
reservoir_weight[139][72],
reservoir_weight[139][73],
reservoir_weight[139][74],
reservoir_weight[139][75],
reservoir_weight[139][76],
reservoir_weight[139][77],
reservoir_weight[139][78],
reservoir_weight[139][79],
reservoir_weight[139][80],
reservoir_weight[139][81],
reservoir_weight[139][82],
reservoir_weight[139][83],
reservoir_weight[139][84],
reservoir_weight[139][85],
reservoir_weight[139][86],
reservoir_weight[139][87],
reservoir_weight[139][88],
reservoir_weight[139][89],
reservoir_weight[139][90],
reservoir_weight[139][91],
reservoir_weight[139][92],
reservoir_weight[139][93],
reservoir_weight[139][94],
reservoir_weight[139][95],
reservoir_weight[139][96],
reservoir_weight[139][97],
reservoir_weight[139][98],
reservoir_weight[139][99],
reservoir_weight[139][100],
reservoir_weight[139][101],
reservoir_weight[139][102],
reservoir_weight[139][103],
reservoir_weight[139][104],
reservoir_weight[139][105],
reservoir_weight[139][106],
reservoir_weight[139][107],
reservoir_weight[139][108],
reservoir_weight[139][109],
reservoir_weight[139][110],
reservoir_weight[139][111],
reservoir_weight[139][112],
reservoir_weight[139][113],
reservoir_weight[139][114],
reservoir_weight[139][115],
reservoir_weight[139][116],
reservoir_weight[139][117],
reservoir_weight[139][118],
reservoir_weight[139][119],
reservoir_weight[139][120],
reservoir_weight[139][121],
reservoir_weight[139][122],
reservoir_weight[139][123],
reservoir_weight[139][124],
reservoir_weight[139][125],
reservoir_weight[139][126],
reservoir_weight[139][127],
reservoir_weight[139][128],
reservoir_weight[139][129],
reservoir_weight[139][130],
reservoir_weight[139][131],
reservoir_weight[139][132],
reservoir_weight[139][133],
reservoir_weight[139][134],
reservoir_weight[139][135],
reservoir_weight[139][136],
reservoir_weight[139][137],
reservoir_weight[139][138],
reservoir_weight[139][139],
reservoir_weight[139][140],
reservoir_weight[139][141],
reservoir_weight[139][142],
reservoir_weight[139][143],
reservoir_weight[139][144],
reservoir_weight[139][145],
reservoir_weight[139][146],
reservoir_weight[139][147],
reservoir_weight[139][148],
reservoir_weight[139][149],
reservoir_weight[139][150],
reservoir_weight[139][151],
reservoir_weight[139][152],
reservoir_weight[139][153],
reservoir_weight[139][154],
reservoir_weight[139][155],
reservoir_weight[139][156],
reservoir_weight[139][157],
reservoir_weight[139][158],
reservoir_weight[139][159],
reservoir_weight[139][160],
reservoir_weight[139][161],
reservoir_weight[139][162],
reservoir_weight[139][163],
reservoir_weight[139][164],
reservoir_weight[139][165],
reservoir_weight[139][166],
reservoir_weight[139][167],
reservoir_weight[139][168],
reservoir_weight[139][169],
reservoir_weight[139][170],
reservoir_weight[139][171],
reservoir_weight[139][172],
reservoir_weight[139][173],
reservoir_weight[139][174],
reservoir_weight[139][175],
reservoir_weight[139][176],
reservoir_weight[139][177],
reservoir_weight[139][178],
reservoir_weight[139][179],
reservoir_weight[139][180],
reservoir_weight[139][181],
reservoir_weight[139][182],
reservoir_weight[139][183],
reservoir_weight[139][184],
reservoir_weight[139][185],
reservoir_weight[139][186],
reservoir_weight[139][187],
reservoir_weight[139][188],
reservoir_weight[139][189],
reservoir_weight[139][190],
reservoir_weight[139][191],
reservoir_weight[139][192],
reservoir_weight[139][193],
reservoir_weight[139][194],
reservoir_weight[139][195],
reservoir_weight[139][196],
reservoir_weight[139][197],
reservoir_weight[139][198],
reservoir_weight[139][199]
},
{reservoir_weight[140][0],
reservoir_weight[140][1],
reservoir_weight[140][2],
reservoir_weight[140][3],
reservoir_weight[140][4],
reservoir_weight[140][5],
reservoir_weight[140][6],
reservoir_weight[140][7],
reservoir_weight[140][8],
reservoir_weight[140][9],
reservoir_weight[140][10],
reservoir_weight[140][11],
reservoir_weight[140][12],
reservoir_weight[140][13],
reservoir_weight[140][14],
reservoir_weight[140][15],
reservoir_weight[140][16],
reservoir_weight[140][17],
reservoir_weight[140][18],
reservoir_weight[140][19],
reservoir_weight[140][20],
reservoir_weight[140][21],
reservoir_weight[140][22],
reservoir_weight[140][23],
reservoir_weight[140][24],
reservoir_weight[140][25],
reservoir_weight[140][26],
reservoir_weight[140][27],
reservoir_weight[140][28],
reservoir_weight[140][29],
reservoir_weight[140][30],
reservoir_weight[140][31],
reservoir_weight[140][32],
reservoir_weight[140][33],
reservoir_weight[140][34],
reservoir_weight[140][35],
reservoir_weight[140][36],
reservoir_weight[140][37],
reservoir_weight[140][38],
reservoir_weight[140][39],
reservoir_weight[140][40],
reservoir_weight[140][41],
reservoir_weight[140][42],
reservoir_weight[140][43],
reservoir_weight[140][44],
reservoir_weight[140][45],
reservoir_weight[140][46],
reservoir_weight[140][47],
reservoir_weight[140][48],
reservoir_weight[140][49],
reservoir_weight[140][50],
reservoir_weight[140][51],
reservoir_weight[140][52],
reservoir_weight[140][53],
reservoir_weight[140][54],
reservoir_weight[140][55],
reservoir_weight[140][56],
reservoir_weight[140][57],
reservoir_weight[140][58],
reservoir_weight[140][59],
reservoir_weight[140][60],
reservoir_weight[140][61],
reservoir_weight[140][62],
reservoir_weight[140][63],
reservoir_weight[140][64],
reservoir_weight[140][65],
reservoir_weight[140][66],
reservoir_weight[140][67],
reservoir_weight[140][68],
reservoir_weight[140][69],
reservoir_weight[140][70],
reservoir_weight[140][71],
reservoir_weight[140][72],
reservoir_weight[140][73],
reservoir_weight[140][74],
reservoir_weight[140][75],
reservoir_weight[140][76],
reservoir_weight[140][77],
reservoir_weight[140][78],
reservoir_weight[140][79],
reservoir_weight[140][80],
reservoir_weight[140][81],
reservoir_weight[140][82],
reservoir_weight[140][83],
reservoir_weight[140][84],
reservoir_weight[140][85],
reservoir_weight[140][86],
reservoir_weight[140][87],
reservoir_weight[140][88],
reservoir_weight[140][89],
reservoir_weight[140][90],
reservoir_weight[140][91],
reservoir_weight[140][92],
reservoir_weight[140][93],
reservoir_weight[140][94],
reservoir_weight[140][95],
reservoir_weight[140][96],
reservoir_weight[140][97],
reservoir_weight[140][98],
reservoir_weight[140][99],
reservoir_weight[140][100],
reservoir_weight[140][101],
reservoir_weight[140][102],
reservoir_weight[140][103],
reservoir_weight[140][104],
reservoir_weight[140][105],
reservoir_weight[140][106],
reservoir_weight[140][107],
reservoir_weight[140][108],
reservoir_weight[140][109],
reservoir_weight[140][110],
reservoir_weight[140][111],
reservoir_weight[140][112],
reservoir_weight[140][113],
reservoir_weight[140][114],
reservoir_weight[140][115],
reservoir_weight[140][116],
reservoir_weight[140][117],
reservoir_weight[140][118],
reservoir_weight[140][119],
reservoir_weight[140][120],
reservoir_weight[140][121],
reservoir_weight[140][122],
reservoir_weight[140][123],
reservoir_weight[140][124],
reservoir_weight[140][125],
reservoir_weight[140][126],
reservoir_weight[140][127],
reservoir_weight[140][128],
reservoir_weight[140][129],
reservoir_weight[140][130],
reservoir_weight[140][131],
reservoir_weight[140][132],
reservoir_weight[140][133],
reservoir_weight[140][134],
reservoir_weight[140][135],
reservoir_weight[140][136],
reservoir_weight[140][137],
reservoir_weight[140][138],
reservoir_weight[140][139],
reservoir_weight[140][140],
reservoir_weight[140][141],
reservoir_weight[140][142],
reservoir_weight[140][143],
reservoir_weight[140][144],
reservoir_weight[140][145],
reservoir_weight[140][146],
reservoir_weight[140][147],
reservoir_weight[140][148],
reservoir_weight[140][149],
reservoir_weight[140][150],
reservoir_weight[140][151],
reservoir_weight[140][152],
reservoir_weight[140][153],
reservoir_weight[140][154],
reservoir_weight[140][155],
reservoir_weight[140][156],
reservoir_weight[140][157],
reservoir_weight[140][158],
reservoir_weight[140][159],
reservoir_weight[140][160],
reservoir_weight[140][161],
reservoir_weight[140][162],
reservoir_weight[140][163],
reservoir_weight[140][164],
reservoir_weight[140][165],
reservoir_weight[140][166],
reservoir_weight[140][167],
reservoir_weight[140][168],
reservoir_weight[140][169],
reservoir_weight[140][170],
reservoir_weight[140][171],
reservoir_weight[140][172],
reservoir_weight[140][173],
reservoir_weight[140][174],
reservoir_weight[140][175],
reservoir_weight[140][176],
reservoir_weight[140][177],
reservoir_weight[140][178],
reservoir_weight[140][179],
reservoir_weight[140][180],
reservoir_weight[140][181],
reservoir_weight[140][182],
reservoir_weight[140][183],
reservoir_weight[140][184],
reservoir_weight[140][185],
reservoir_weight[140][186],
reservoir_weight[140][187],
reservoir_weight[140][188],
reservoir_weight[140][189],
reservoir_weight[140][190],
reservoir_weight[140][191],
reservoir_weight[140][192],
reservoir_weight[140][193],
reservoir_weight[140][194],
reservoir_weight[140][195],
reservoir_weight[140][196],
reservoir_weight[140][197],
reservoir_weight[140][198],
reservoir_weight[140][199]
},
{reservoir_weight[141][0],
reservoir_weight[141][1],
reservoir_weight[141][2],
reservoir_weight[141][3],
reservoir_weight[141][4],
reservoir_weight[141][5],
reservoir_weight[141][6],
reservoir_weight[141][7],
reservoir_weight[141][8],
reservoir_weight[141][9],
reservoir_weight[141][10],
reservoir_weight[141][11],
reservoir_weight[141][12],
reservoir_weight[141][13],
reservoir_weight[141][14],
reservoir_weight[141][15],
reservoir_weight[141][16],
reservoir_weight[141][17],
reservoir_weight[141][18],
reservoir_weight[141][19],
reservoir_weight[141][20],
reservoir_weight[141][21],
reservoir_weight[141][22],
reservoir_weight[141][23],
reservoir_weight[141][24],
reservoir_weight[141][25],
reservoir_weight[141][26],
reservoir_weight[141][27],
reservoir_weight[141][28],
reservoir_weight[141][29],
reservoir_weight[141][30],
reservoir_weight[141][31],
reservoir_weight[141][32],
reservoir_weight[141][33],
reservoir_weight[141][34],
reservoir_weight[141][35],
reservoir_weight[141][36],
reservoir_weight[141][37],
reservoir_weight[141][38],
reservoir_weight[141][39],
reservoir_weight[141][40],
reservoir_weight[141][41],
reservoir_weight[141][42],
reservoir_weight[141][43],
reservoir_weight[141][44],
reservoir_weight[141][45],
reservoir_weight[141][46],
reservoir_weight[141][47],
reservoir_weight[141][48],
reservoir_weight[141][49],
reservoir_weight[141][50],
reservoir_weight[141][51],
reservoir_weight[141][52],
reservoir_weight[141][53],
reservoir_weight[141][54],
reservoir_weight[141][55],
reservoir_weight[141][56],
reservoir_weight[141][57],
reservoir_weight[141][58],
reservoir_weight[141][59],
reservoir_weight[141][60],
reservoir_weight[141][61],
reservoir_weight[141][62],
reservoir_weight[141][63],
reservoir_weight[141][64],
reservoir_weight[141][65],
reservoir_weight[141][66],
reservoir_weight[141][67],
reservoir_weight[141][68],
reservoir_weight[141][69],
reservoir_weight[141][70],
reservoir_weight[141][71],
reservoir_weight[141][72],
reservoir_weight[141][73],
reservoir_weight[141][74],
reservoir_weight[141][75],
reservoir_weight[141][76],
reservoir_weight[141][77],
reservoir_weight[141][78],
reservoir_weight[141][79],
reservoir_weight[141][80],
reservoir_weight[141][81],
reservoir_weight[141][82],
reservoir_weight[141][83],
reservoir_weight[141][84],
reservoir_weight[141][85],
reservoir_weight[141][86],
reservoir_weight[141][87],
reservoir_weight[141][88],
reservoir_weight[141][89],
reservoir_weight[141][90],
reservoir_weight[141][91],
reservoir_weight[141][92],
reservoir_weight[141][93],
reservoir_weight[141][94],
reservoir_weight[141][95],
reservoir_weight[141][96],
reservoir_weight[141][97],
reservoir_weight[141][98],
reservoir_weight[141][99],
reservoir_weight[141][100],
reservoir_weight[141][101],
reservoir_weight[141][102],
reservoir_weight[141][103],
reservoir_weight[141][104],
reservoir_weight[141][105],
reservoir_weight[141][106],
reservoir_weight[141][107],
reservoir_weight[141][108],
reservoir_weight[141][109],
reservoir_weight[141][110],
reservoir_weight[141][111],
reservoir_weight[141][112],
reservoir_weight[141][113],
reservoir_weight[141][114],
reservoir_weight[141][115],
reservoir_weight[141][116],
reservoir_weight[141][117],
reservoir_weight[141][118],
reservoir_weight[141][119],
reservoir_weight[141][120],
reservoir_weight[141][121],
reservoir_weight[141][122],
reservoir_weight[141][123],
reservoir_weight[141][124],
reservoir_weight[141][125],
reservoir_weight[141][126],
reservoir_weight[141][127],
reservoir_weight[141][128],
reservoir_weight[141][129],
reservoir_weight[141][130],
reservoir_weight[141][131],
reservoir_weight[141][132],
reservoir_weight[141][133],
reservoir_weight[141][134],
reservoir_weight[141][135],
reservoir_weight[141][136],
reservoir_weight[141][137],
reservoir_weight[141][138],
reservoir_weight[141][139],
reservoir_weight[141][140],
reservoir_weight[141][141],
reservoir_weight[141][142],
reservoir_weight[141][143],
reservoir_weight[141][144],
reservoir_weight[141][145],
reservoir_weight[141][146],
reservoir_weight[141][147],
reservoir_weight[141][148],
reservoir_weight[141][149],
reservoir_weight[141][150],
reservoir_weight[141][151],
reservoir_weight[141][152],
reservoir_weight[141][153],
reservoir_weight[141][154],
reservoir_weight[141][155],
reservoir_weight[141][156],
reservoir_weight[141][157],
reservoir_weight[141][158],
reservoir_weight[141][159],
reservoir_weight[141][160],
reservoir_weight[141][161],
reservoir_weight[141][162],
reservoir_weight[141][163],
reservoir_weight[141][164],
reservoir_weight[141][165],
reservoir_weight[141][166],
reservoir_weight[141][167],
reservoir_weight[141][168],
reservoir_weight[141][169],
reservoir_weight[141][170],
reservoir_weight[141][171],
reservoir_weight[141][172],
reservoir_weight[141][173],
reservoir_weight[141][174],
reservoir_weight[141][175],
reservoir_weight[141][176],
reservoir_weight[141][177],
reservoir_weight[141][178],
reservoir_weight[141][179],
reservoir_weight[141][180],
reservoir_weight[141][181],
reservoir_weight[141][182],
reservoir_weight[141][183],
reservoir_weight[141][184],
reservoir_weight[141][185],
reservoir_weight[141][186],
reservoir_weight[141][187],
reservoir_weight[141][188],
reservoir_weight[141][189],
reservoir_weight[141][190],
reservoir_weight[141][191],
reservoir_weight[141][192],
reservoir_weight[141][193],
reservoir_weight[141][194],
reservoir_weight[141][195],
reservoir_weight[141][196],
reservoir_weight[141][197],
reservoir_weight[141][198],
reservoir_weight[141][199]
},
{reservoir_weight[142][0],
reservoir_weight[142][1],
reservoir_weight[142][2],
reservoir_weight[142][3],
reservoir_weight[142][4],
reservoir_weight[142][5],
reservoir_weight[142][6],
reservoir_weight[142][7],
reservoir_weight[142][8],
reservoir_weight[142][9],
reservoir_weight[142][10],
reservoir_weight[142][11],
reservoir_weight[142][12],
reservoir_weight[142][13],
reservoir_weight[142][14],
reservoir_weight[142][15],
reservoir_weight[142][16],
reservoir_weight[142][17],
reservoir_weight[142][18],
reservoir_weight[142][19],
reservoir_weight[142][20],
reservoir_weight[142][21],
reservoir_weight[142][22],
reservoir_weight[142][23],
reservoir_weight[142][24],
reservoir_weight[142][25],
reservoir_weight[142][26],
reservoir_weight[142][27],
reservoir_weight[142][28],
reservoir_weight[142][29],
reservoir_weight[142][30],
reservoir_weight[142][31],
reservoir_weight[142][32],
reservoir_weight[142][33],
reservoir_weight[142][34],
reservoir_weight[142][35],
reservoir_weight[142][36],
reservoir_weight[142][37],
reservoir_weight[142][38],
reservoir_weight[142][39],
reservoir_weight[142][40],
reservoir_weight[142][41],
reservoir_weight[142][42],
reservoir_weight[142][43],
reservoir_weight[142][44],
reservoir_weight[142][45],
reservoir_weight[142][46],
reservoir_weight[142][47],
reservoir_weight[142][48],
reservoir_weight[142][49],
reservoir_weight[142][50],
reservoir_weight[142][51],
reservoir_weight[142][52],
reservoir_weight[142][53],
reservoir_weight[142][54],
reservoir_weight[142][55],
reservoir_weight[142][56],
reservoir_weight[142][57],
reservoir_weight[142][58],
reservoir_weight[142][59],
reservoir_weight[142][60],
reservoir_weight[142][61],
reservoir_weight[142][62],
reservoir_weight[142][63],
reservoir_weight[142][64],
reservoir_weight[142][65],
reservoir_weight[142][66],
reservoir_weight[142][67],
reservoir_weight[142][68],
reservoir_weight[142][69],
reservoir_weight[142][70],
reservoir_weight[142][71],
reservoir_weight[142][72],
reservoir_weight[142][73],
reservoir_weight[142][74],
reservoir_weight[142][75],
reservoir_weight[142][76],
reservoir_weight[142][77],
reservoir_weight[142][78],
reservoir_weight[142][79],
reservoir_weight[142][80],
reservoir_weight[142][81],
reservoir_weight[142][82],
reservoir_weight[142][83],
reservoir_weight[142][84],
reservoir_weight[142][85],
reservoir_weight[142][86],
reservoir_weight[142][87],
reservoir_weight[142][88],
reservoir_weight[142][89],
reservoir_weight[142][90],
reservoir_weight[142][91],
reservoir_weight[142][92],
reservoir_weight[142][93],
reservoir_weight[142][94],
reservoir_weight[142][95],
reservoir_weight[142][96],
reservoir_weight[142][97],
reservoir_weight[142][98],
reservoir_weight[142][99],
reservoir_weight[142][100],
reservoir_weight[142][101],
reservoir_weight[142][102],
reservoir_weight[142][103],
reservoir_weight[142][104],
reservoir_weight[142][105],
reservoir_weight[142][106],
reservoir_weight[142][107],
reservoir_weight[142][108],
reservoir_weight[142][109],
reservoir_weight[142][110],
reservoir_weight[142][111],
reservoir_weight[142][112],
reservoir_weight[142][113],
reservoir_weight[142][114],
reservoir_weight[142][115],
reservoir_weight[142][116],
reservoir_weight[142][117],
reservoir_weight[142][118],
reservoir_weight[142][119],
reservoir_weight[142][120],
reservoir_weight[142][121],
reservoir_weight[142][122],
reservoir_weight[142][123],
reservoir_weight[142][124],
reservoir_weight[142][125],
reservoir_weight[142][126],
reservoir_weight[142][127],
reservoir_weight[142][128],
reservoir_weight[142][129],
reservoir_weight[142][130],
reservoir_weight[142][131],
reservoir_weight[142][132],
reservoir_weight[142][133],
reservoir_weight[142][134],
reservoir_weight[142][135],
reservoir_weight[142][136],
reservoir_weight[142][137],
reservoir_weight[142][138],
reservoir_weight[142][139],
reservoir_weight[142][140],
reservoir_weight[142][141],
reservoir_weight[142][142],
reservoir_weight[142][143],
reservoir_weight[142][144],
reservoir_weight[142][145],
reservoir_weight[142][146],
reservoir_weight[142][147],
reservoir_weight[142][148],
reservoir_weight[142][149],
reservoir_weight[142][150],
reservoir_weight[142][151],
reservoir_weight[142][152],
reservoir_weight[142][153],
reservoir_weight[142][154],
reservoir_weight[142][155],
reservoir_weight[142][156],
reservoir_weight[142][157],
reservoir_weight[142][158],
reservoir_weight[142][159],
reservoir_weight[142][160],
reservoir_weight[142][161],
reservoir_weight[142][162],
reservoir_weight[142][163],
reservoir_weight[142][164],
reservoir_weight[142][165],
reservoir_weight[142][166],
reservoir_weight[142][167],
reservoir_weight[142][168],
reservoir_weight[142][169],
reservoir_weight[142][170],
reservoir_weight[142][171],
reservoir_weight[142][172],
reservoir_weight[142][173],
reservoir_weight[142][174],
reservoir_weight[142][175],
reservoir_weight[142][176],
reservoir_weight[142][177],
reservoir_weight[142][178],
reservoir_weight[142][179],
reservoir_weight[142][180],
reservoir_weight[142][181],
reservoir_weight[142][182],
reservoir_weight[142][183],
reservoir_weight[142][184],
reservoir_weight[142][185],
reservoir_weight[142][186],
reservoir_weight[142][187],
reservoir_weight[142][188],
reservoir_weight[142][189],
reservoir_weight[142][190],
reservoir_weight[142][191],
reservoir_weight[142][192],
reservoir_weight[142][193],
reservoir_weight[142][194],
reservoir_weight[142][195],
reservoir_weight[142][196],
reservoir_weight[142][197],
reservoir_weight[142][198],
reservoir_weight[142][199]
},
{reservoir_weight[143][0],
reservoir_weight[143][1],
reservoir_weight[143][2],
reservoir_weight[143][3],
reservoir_weight[143][4],
reservoir_weight[143][5],
reservoir_weight[143][6],
reservoir_weight[143][7],
reservoir_weight[143][8],
reservoir_weight[143][9],
reservoir_weight[143][10],
reservoir_weight[143][11],
reservoir_weight[143][12],
reservoir_weight[143][13],
reservoir_weight[143][14],
reservoir_weight[143][15],
reservoir_weight[143][16],
reservoir_weight[143][17],
reservoir_weight[143][18],
reservoir_weight[143][19],
reservoir_weight[143][20],
reservoir_weight[143][21],
reservoir_weight[143][22],
reservoir_weight[143][23],
reservoir_weight[143][24],
reservoir_weight[143][25],
reservoir_weight[143][26],
reservoir_weight[143][27],
reservoir_weight[143][28],
reservoir_weight[143][29],
reservoir_weight[143][30],
reservoir_weight[143][31],
reservoir_weight[143][32],
reservoir_weight[143][33],
reservoir_weight[143][34],
reservoir_weight[143][35],
reservoir_weight[143][36],
reservoir_weight[143][37],
reservoir_weight[143][38],
reservoir_weight[143][39],
reservoir_weight[143][40],
reservoir_weight[143][41],
reservoir_weight[143][42],
reservoir_weight[143][43],
reservoir_weight[143][44],
reservoir_weight[143][45],
reservoir_weight[143][46],
reservoir_weight[143][47],
reservoir_weight[143][48],
reservoir_weight[143][49],
reservoir_weight[143][50],
reservoir_weight[143][51],
reservoir_weight[143][52],
reservoir_weight[143][53],
reservoir_weight[143][54],
reservoir_weight[143][55],
reservoir_weight[143][56],
reservoir_weight[143][57],
reservoir_weight[143][58],
reservoir_weight[143][59],
reservoir_weight[143][60],
reservoir_weight[143][61],
reservoir_weight[143][62],
reservoir_weight[143][63],
reservoir_weight[143][64],
reservoir_weight[143][65],
reservoir_weight[143][66],
reservoir_weight[143][67],
reservoir_weight[143][68],
reservoir_weight[143][69],
reservoir_weight[143][70],
reservoir_weight[143][71],
reservoir_weight[143][72],
reservoir_weight[143][73],
reservoir_weight[143][74],
reservoir_weight[143][75],
reservoir_weight[143][76],
reservoir_weight[143][77],
reservoir_weight[143][78],
reservoir_weight[143][79],
reservoir_weight[143][80],
reservoir_weight[143][81],
reservoir_weight[143][82],
reservoir_weight[143][83],
reservoir_weight[143][84],
reservoir_weight[143][85],
reservoir_weight[143][86],
reservoir_weight[143][87],
reservoir_weight[143][88],
reservoir_weight[143][89],
reservoir_weight[143][90],
reservoir_weight[143][91],
reservoir_weight[143][92],
reservoir_weight[143][93],
reservoir_weight[143][94],
reservoir_weight[143][95],
reservoir_weight[143][96],
reservoir_weight[143][97],
reservoir_weight[143][98],
reservoir_weight[143][99],
reservoir_weight[143][100],
reservoir_weight[143][101],
reservoir_weight[143][102],
reservoir_weight[143][103],
reservoir_weight[143][104],
reservoir_weight[143][105],
reservoir_weight[143][106],
reservoir_weight[143][107],
reservoir_weight[143][108],
reservoir_weight[143][109],
reservoir_weight[143][110],
reservoir_weight[143][111],
reservoir_weight[143][112],
reservoir_weight[143][113],
reservoir_weight[143][114],
reservoir_weight[143][115],
reservoir_weight[143][116],
reservoir_weight[143][117],
reservoir_weight[143][118],
reservoir_weight[143][119],
reservoir_weight[143][120],
reservoir_weight[143][121],
reservoir_weight[143][122],
reservoir_weight[143][123],
reservoir_weight[143][124],
reservoir_weight[143][125],
reservoir_weight[143][126],
reservoir_weight[143][127],
reservoir_weight[143][128],
reservoir_weight[143][129],
reservoir_weight[143][130],
reservoir_weight[143][131],
reservoir_weight[143][132],
reservoir_weight[143][133],
reservoir_weight[143][134],
reservoir_weight[143][135],
reservoir_weight[143][136],
reservoir_weight[143][137],
reservoir_weight[143][138],
reservoir_weight[143][139],
reservoir_weight[143][140],
reservoir_weight[143][141],
reservoir_weight[143][142],
reservoir_weight[143][143],
reservoir_weight[143][144],
reservoir_weight[143][145],
reservoir_weight[143][146],
reservoir_weight[143][147],
reservoir_weight[143][148],
reservoir_weight[143][149],
reservoir_weight[143][150],
reservoir_weight[143][151],
reservoir_weight[143][152],
reservoir_weight[143][153],
reservoir_weight[143][154],
reservoir_weight[143][155],
reservoir_weight[143][156],
reservoir_weight[143][157],
reservoir_weight[143][158],
reservoir_weight[143][159],
reservoir_weight[143][160],
reservoir_weight[143][161],
reservoir_weight[143][162],
reservoir_weight[143][163],
reservoir_weight[143][164],
reservoir_weight[143][165],
reservoir_weight[143][166],
reservoir_weight[143][167],
reservoir_weight[143][168],
reservoir_weight[143][169],
reservoir_weight[143][170],
reservoir_weight[143][171],
reservoir_weight[143][172],
reservoir_weight[143][173],
reservoir_weight[143][174],
reservoir_weight[143][175],
reservoir_weight[143][176],
reservoir_weight[143][177],
reservoir_weight[143][178],
reservoir_weight[143][179],
reservoir_weight[143][180],
reservoir_weight[143][181],
reservoir_weight[143][182],
reservoir_weight[143][183],
reservoir_weight[143][184],
reservoir_weight[143][185],
reservoir_weight[143][186],
reservoir_weight[143][187],
reservoir_weight[143][188],
reservoir_weight[143][189],
reservoir_weight[143][190],
reservoir_weight[143][191],
reservoir_weight[143][192],
reservoir_weight[143][193],
reservoir_weight[143][194],
reservoir_weight[143][195],
reservoir_weight[143][196],
reservoir_weight[143][197],
reservoir_weight[143][198],
reservoir_weight[143][199]
},
{reservoir_weight[144][0],
reservoir_weight[144][1],
reservoir_weight[144][2],
reservoir_weight[144][3],
reservoir_weight[144][4],
reservoir_weight[144][5],
reservoir_weight[144][6],
reservoir_weight[144][7],
reservoir_weight[144][8],
reservoir_weight[144][9],
reservoir_weight[144][10],
reservoir_weight[144][11],
reservoir_weight[144][12],
reservoir_weight[144][13],
reservoir_weight[144][14],
reservoir_weight[144][15],
reservoir_weight[144][16],
reservoir_weight[144][17],
reservoir_weight[144][18],
reservoir_weight[144][19],
reservoir_weight[144][20],
reservoir_weight[144][21],
reservoir_weight[144][22],
reservoir_weight[144][23],
reservoir_weight[144][24],
reservoir_weight[144][25],
reservoir_weight[144][26],
reservoir_weight[144][27],
reservoir_weight[144][28],
reservoir_weight[144][29],
reservoir_weight[144][30],
reservoir_weight[144][31],
reservoir_weight[144][32],
reservoir_weight[144][33],
reservoir_weight[144][34],
reservoir_weight[144][35],
reservoir_weight[144][36],
reservoir_weight[144][37],
reservoir_weight[144][38],
reservoir_weight[144][39],
reservoir_weight[144][40],
reservoir_weight[144][41],
reservoir_weight[144][42],
reservoir_weight[144][43],
reservoir_weight[144][44],
reservoir_weight[144][45],
reservoir_weight[144][46],
reservoir_weight[144][47],
reservoir_weight[144][48],
reservoir_weight[144][49],
reservoir_weight[144][50],
reservoir_weight[144][51],
reservoir_weight[144][52],
reservoir_weight[144][53],
reservoir_weight[144][54],
reservoir_weight[144][55],
reservoir_weight[144][56],
reservoir_weight[144][57],
reservoir_weight[144][58],
reservoir_weight[144][59],
reservoir_weight[144][60],
reservoir_weight[144][61],
reservoir_weight[144][62],
reservoir_weight[144][63],
reservoir_weight[144][64],
reservoir_weight[144][65],
reservoir_weight[144][66],
reservoir_weight[144][67],
reservoir_weight[144][68],
reservoir_weight[144][69],
reservoir_weight[144][70],
reservoir_weight[144][71],
reservoir_weight[144][72],
reservoir_weight[144][73],
reservoir_weight[144][74],
reservoir_weight[144][75],
reservoir_weight[144][76],
reservoir_weight[144][77],
reservoir_weight[144][78],
reservoir_weight[144][79],
reservoir_weight[144][80],
reservoir_weight[144][81],
reservoir_weight[144][82],
reservoir_weight[144][83],
reservoir_weight[144][84],
reservoir_weight[144][85],
reservoir_weight[144][86],
reservoir_weight[144][87],
reservoir_weight[144][88],
reservoir_weight[144][89],
reservoir_weight[144][90],
reservoir_weight[144][91],
reservoir_weight[144][92],
reservoir_weight[144][93],
reservoir_weight[144][94],
reservoir_weight[144][95],
reservoir_weight[144][96],
reservoir_weight[144][97],
reservoir_weight[144][98],
reservoir_weight[144][99],
reservoir_weight[144][100],
reservoir_weight[144][101],
reservoir_weight[144][102],
reservoir_weight[144][103],
reservoir_weight[144][104],
reservoir_weight[144][105],
reservoir_weight[144][106],
reservoir_weight[144][107],
reservoir_weight[144][108],
reservoir_weight[144][109],
reservoir_weight[144][110],
reservoir_weight[144][111],
reservoir_weight[144][112],
reservoir_weight[144][113],
reservoir_weight[144][114],
reservoir_weight[144][115],
reservoir_weight[144][116],
reservoir_weight[144][117],
reservoir_weight[144][118],
reservoir_weight[144][119],
reservoir_weight[144][120],
reservoir_weight[144][121],
reservoir_weight[144][122],
reservoir_weight[144][123],
reservoir_weight[144][124],
reservoir_weight[144][125],
reservoir_weight[144][126],
reservoir_weight[144][127],
reservoir_weight[144][128],
reservoir_weight[144][129],
reservoir_weight[144][130],
reservoir_weight[144][131],
reservoir_weight[144][132],
reservoir_weight[144][133],
reservoir_weight[144][134],
reservoir_weight[144][135],
reservoir_weight[144][136],
reservoir_weight[144][137],
reservoir_weight[144][138],
reservoir_weight[144][139],
reservoir_weight[144][140],
reservoir_weight[144][141],
reservoir_weight[144][142],
reservoir_weight[144][143],
reservoir_weight[144][144],
reservoir_weight[144][145],
reservoir_weight[144][146],
reservoir_weight[144][147],
reservoir_weight[144][148],
reservoir_weight[144][149],
reservoir_weight[144][150],
reservoir_weight[144][151],
reservoir_weight[144][152],
reservoir_weight[144][153],
reservoir_weight[144][154],
reservoir_weight[144][155],
reservoir_weight[144][156],
reservoir_weight[144][157],
reservoir_weight[144][158],
reservoir_weight[144][159],
reservoir_weight[144][160],
reservoir_weight[144][161],
reservoir_weight[144][162],
reservoir_weight[144][163],
reservoir_weight[144][164],
reservoir_weight[144][165],
reservoir_weight[144][166],
reservoir_weight[144][167],
reservoir_weight[144][168],
reservoir_weight[144][169],
reservoir_weight[144][170],
reservoir_weight[144][171],
reservoir_weight[144][172],
reservoir_weight[144][173],
reservoir_weight[144][174],
reservoir_weight[144][175],
reservoir_weight[144][176],
reservoir_weight[144][177],
reservoir_weight[144][178],
reservoir_weight[144][179],
reservoir_weight[144][180],
reservoir_weight[144][181],
reservoir_weight[144][182],
reservoir_weight[144][183],
reservoir_weight[144][184],
reservoir_weight[144][185],
reservoir_weight[144][186],
reservoir_weight[144][187],
reservoir_weight[144][188],
reservoir_weight[144][189],
reservoir_weight[144][190],
reservoir_weight[144][191],
reservoir_weight[144][192],
reservoir_weight[144][193],
reservoir_weight[144][194],
reservoir_weight[144][195],
reservoir_weight[144][196],
reservoir_weight[144][197],
reservoir_weight[144][198],
reservoir_weight[144][199]
},
{reservoir_weight[145][0],
reservoir_weight[145][1],
reservoir_weight[145][2],
reservoir_weight[145][3],
reservoir_weight[145][4],
reservoir_weight[145][5],
reservoir_weight[145][6],
reservoir_weight[145][7],
reservoir_weight[145][8],
reservoir_weight[145][9],
reservoir_weight[145][10],
reservoir_weight[145][11],
reservoir_weight[145][12],
reservoir_weight[145][13],
reservoir_weight[145][14],
reservoir_weight[145][15],
reservoir_weight[145][16],
reservoir_weight[145][17],
reservoir_weight[145][18],
reservoir_weight[145][19],
reservoir_weight[145][20],
reservoir_weight[145][21],
reservoir_weight[145][22],
reservoir_weight[145][23],
reservoir_weight[145][24],
reservoir_weight[145][25],
reservoir_weight[145][26],
reservoir_weight[145][27],
reservoir_weight[145][28],
reservoir_weight[145][29],
reservoir_weight[145][30],
reservoir_weight[145][31],
reservoir_weight[145][32],
reservoir_weight[145][33],
reservoir_weight[145][34],
reservoir_weight[145][35],
reservoir_weight[145][36],
reservoir_weight[145][37],
reservoir_weight[145][38],
reservoir_weight[145][39],
reservoir_weight[145][40],
reservoir_weight[145][41],
reservoir_weight[145][42],
reservoir_weight[145][43],
reservoir_weight[145][44],
reservoir_weight[145][45],
reservoir_weight[145][46],
reservoir_weight[145][47],
reservoir_weight[145][48],
reservoir_weight[145][49],
reservoir_weight[145][50],
reservoir_weight[145][51],
reservoir_weight[145][52],
reservoir_weight[145][53],
reservoir_weight[145][54],
reservoir_weight[145][55],
reservoir_weight[145][56],
reservoir_weight[145][57],
reservoir_weight[145][58],
reservoir_weight[145][59],
reservoir_weight[145][60],
reservoir_weight[145][61],
reservoir_weight[145][62],
reservoir_weight[145][63],
reservoir_weight[145][64],
reservoir_weight[145][65],
reservoir_weight[145][66],
reservoir_weight[145][67],
reservoir_weight[145][68],
reservoir_weight[145][69],
reservoir_weight[145][70],
reservoir_weight[145][71],
reservoir_weight[145][72],
reservoir_weight[145][73],
reservoir_weight[145][74],
reservoir_weight[145][75],
reservoir_weight[145][76],
reservoir_weight[145][77],
reservoir_weight[145][78],
reservoir_weight[145][79],
reservoir_weight[145][80],
reservoir_weight[145][81],
reservoir_weight[145][82],
reservoir_weight[145][83],
reservoir_weight[145][84],
reservoir_weight[145][85],
reservoir_weight[145][86],
reservoir_weight[145][87],
reservoir_weight[145][88],
reservoir_weight[145][89],
reservoir_weight[145][90],
reservoir_weight[145][91],
reservoir_weight[145][92],
reservoir_weight[145][93],
reservoir_weight[145][94],
reservoir_weight[145][95],
reservoir_weight[145][96],
reservoir_weight[145][97],
reservoir_weight[145][98],
reservoir_weight[145][99],
reservoir_weight[145][100],
reservoir_weight[145][101],
reservoir_weight[145][102],
reservoir_weight[145][103],
reservoir_weight[145][104],
reservoir_weight[145][105],
reservoir_weight[145][106],
reservoir_weight[145][107],
reservoir_weight[145][108],
reservoir_weight[145][109],
reservoir_weight[145][110],
reservoir_weight[145][111],
reservoir_weight[145][112],
reservoir_weight[145][113],
reservoir_weight[145][114],
reservoir_weight[145][115],
reservoir_weight[145][116],
reservoir_weight[145][117],
reservoir_weight[145][118],
reservoir_weight[145][119],
reservoir_weight[145][120],
reservoir_weight[145][121],
reservoir_weight[145][122],
reservoir_weight[145][123],
reservoir_weight[145][124],
reservoir_weight[145][125],
reservoir_weight[145][126],
reservoir_weight[145][127],
reservoir_weight[145][128],
reservoir_weight[145][129],
reservoir_weight[145][130],
reservoir_weight[145][131],
reservoir_weight[145][132],
reservoir_weight[145][133],
reservoir_weight[145][134],
reservoir_weight[145][135],
reservoir_weight[145][136],
reservoir_weight[145][137],
reservoir_weight[145][138],
reservoir_weight[145][139],
reservoir_weight[145][140],
reservoir_weight[145][141],
reservoir_weight[145][142],
reservoir_weight[145][143],
reservoir_weight[145][144],
reservoir_weight[145][145],
reservoir_weight[145][146],
reservoir_weight[145][147],
reservoir_weight[145][148],
reservoir_weight[145][149],
reservoir_weight[145][150],
reservoir_weight[145][151],
reservoir_weight[145][152],
reservoir_weight[145][153],
reservoir_weight[145][154],
reservoir_weight[145][155],
reservoir_weight[145][156],
reservoir_weight[145][157],
reservoir_weight[145][158],
reservoir_weight[145][159],
reservoir_weight[145][160],
reservoir_weight[145][161],
reservoir_weight[145][162],
reservoir_weight[145][163],
reservoir_weight[145][164],
reservoir_weight[145][165],
reservoir_weight[145][166],
reservoir_weight[145][167],
reservoir_weight[145][168],
reservoir_weight[145][169],
reservoir_weight[145][170],
reservoir_weight[145][171],
reservoir_weight[145][172],
reservoir_weight[145][173],
reservoir_weight[145][174],
reservoir_weight[145][175],
reservoir_weight[145][176],
reservoir_weight[145][177],
reservoir_weight[145][178],
reservoir_weight[145][179],
reservoir_weight[145][180],
reservoir_weight[145][181],
reservoir_weight[145][182],
reservoir_weight[145][183],
reservoir_weight[145][184],
reservoir_weight[145][185],
reservoir_weight[145][186],
reservoir_weight[145][187],
reservoir_weight[145][188],
reservoir_weight[145][189],
reservoir_weight[145][190],
reservoir_weight[145][191],
reservoir_weight[145][192],
reservoir_weight[145][193],
reservoir_weight[145][194],
reservoir_weight[145][195],
reservoir_weight[145][196],
reservoir_weight[145][197],
reservoir_weight[145][198],
reservoir_weight[145][199]
},
{reservoir_weight[146][0],
reservoir_weight[146][1],
reservoir_weight[146][2],
reservoir_weight[146][3],
reservoir_weight[146][4],
reservoir_weight[146][5],
reservoir_weight[146][6],
reservoir_weight[146][7],
reservoir_weight[146][8],
reservoir_weight[146][9],
reservoir_weight[146][10],
reservoir_weight[146][11],
reservoir_weight[146][12],
reservoir_weight[146][13],
reservoir_weight[146][14],
reservoir_weight[146][15],
reservoir_weight[146][16],
reservoir_weight[146][17],
reservoir_weight[146][18],
reservoir_weight[146][19],
reservoir_weight[146][20],
reservoir_weight[146][21],
reservoir_weight[146][22],
reservoir_weight[146][23],
reservoir_weight[146][24],
reservoir_weight[146][25],
reservoir_weight[146][26],
reservoir_weight[146][27],
reservoir_weight[146][28],
reservoir_weight[146][29],
reservoir_weight[146][30],
reservoir_weight[146][31],
reservoir_weight[146][32],
reservoir_weight[146][33],
reservoir_weight[146][34],
reservoir_weight[146][35],
reservoir_weight[146][36],
reservoir_weight[146][37],
reservoir_weight[146][38],
reservoir_weight[146][39],
reservoir_weight[146][40],
reservoir_weight[146][41],
reservoir_weight[146][42],
reservoir_weight[146][43],
reservoir_weight[146][44],
reservoir_weight[146][45],
reservoir_weight[146][46],
reservoir_weight[146][47],
reservoir_weight[146][48],
reservoir_weight[146][49],
reservoir_weight[146][50],
reservoir_weight[146][51],
reservoir_weight[146][52],
reservoir_weight[146][53],
reservoir_weight[146][54],
reservoir_weight[146][55],
reservoir_weight[146][56],
reservoir_weight[146][57],
reservoir_weight[146][58],
reservoir_weight[146][59],
reservoir_weight[146][60],
reservoir_weight[146][61],
reservoir_weight[146][62],
reservoir_weight[146][63],
reservoir_weight[146][64],
reservoir_weight[146][65],
reservoir_weight[146][66],
reservoir_weight[146][67],
reservoir_weight[146][68],
reservoir_weight[146][69],
reservoir_weight[146][70],
reservoir_weight[146][71],
reservoir_weight[146][72],
reservoir_weight[146][73],
reservoir_weight[146][74],
reservoir_weight[146][75],
reservoir_weight[146][76],
reservoir_weight[146][77],
reservoir_weight[146][78],
reservoir_weight[146][79],
reservoir_weight[146][80],
reservoir_weight[146][81],
reservoir_weight[146][82],
reservoir_weight[146][83],
reservoir_weight[146][84],
reservoir_weight[146][85],
reservoir_weight[146][86],
reservoir_weight[146][87],
reservoir_weight[146][88],
reservoir_weight[146][89],
reservoir_weight[146][90],
reservoir_weight[146][91],
reservoir_weight[146][92],
reservoir_weight[146][93],
reservoir_weight[146][94],
reservoir_weight[146][95],
reservoir_weight[146][96],
reservoir_weight[146][97],
reservoir_weight[146][98],
reservoir_weight[146][99],
reservoir_weight[146][100],
reservoir_weight[146][101],
reservoir_weight[146][102],
reservoir_weight[146][103],
reservoir_weight[146][104],
reservoir_weight[146][105],
reservoir_weight[146][106],
reservoir_weight[146][107],
reservoir_weight[146][108],
reservoir_weight[146][109],
reservoir_weight[146][110],
reservoir_weight[146][111],
reservoir_weight[146][112],
reservoir_weight[146][113],
reservoir_weight[146][114],
reservoir_weight[146][115],
reservoir_weight[146][116],
reservoir_weight[146][117],
reservoir_weight[146][118],
reservoir_weight[146][119],
reservoir_weight[146][120],
reservoir_weight[146][121],
reservoir_weight[146][122],
reservoir_weight[146][123],
reservoir_weight[146][124],
reservoir_weight[146][125],
reservoir_weight[146][126],
reservoir_weight[146][127],
reservoir_weight[146][128],
reservoir_weight[146][129],
reservoir_weight[146][130],
reservoir_weight[146][131],
reservoir_weight[146][132],
reservoir_weight[146][133],
reservoir_weight[146][134],
reservoir_weight[146][135],
reservoir_weight[146][136],
reservoir_weight[146][137],
reservoir_weight[146][138],
reservoir_weight[146][139],
reservoir_weight[146][140],
reservoir_weight[146][141],
reservoir_weight[146][142],
reservoir_weight[146][143],
reservoir_weight[146][144],
reservoir_weight[146][145],
reservoir_weight[146][146],
reservoir_weight[146][147],
reservoir_weight[146][148],
reservoir_weight[146][149],
reservoir_weight[146][150],
reservoir_weight[146][151],
reservoir_weight[146][152],
reservoir_weight[146][153],
reservoir_weight[146][154],
reservoir_weight[146][155],
reservoir_weight[146][156],
reservoir_weight[146][157],
reservoir_weight[146][158],
reservoir_weight[146][159],
reservoir_weight[146][160],
reservoir_weight[146][161],
reservoir_weight[146][162],
reservoir_weight[146][163],
reservoir_weight[146][164],
reservoir_weight[146][165],
reservoir_weight[146][166],
reservoir_weight[146][167],
reservoir_weight[146][168],
reservoir_weight[146][169],
reservoir_weight[146][170],
reservoir_weight[146][171],
reservoir_weight[146][172],
reservoir_weight[146][173],
reservoir_weight[146][174],
reservoir_weight[146][175],
reservoir_weight[146][176],
reservoir_weight[146][177],
reservoir_weight[146][178],
reservoir_weight[146][179],
reservoir_weight[146][180],
reservoir_weight[146][181],
reservoir_weight[146][182],
reservoir_weight[146][183],
reservoir_weight[146][184],
reservoir_weight[146][185],
reservoir_weight[146][186],
reservoir_weight[146][187],
reservoir_weight[146][188],
reservoir_weight[146][189],
reservoir_weight[146][190],
reservoir_weight[146][191],
reservoir_weight[146][192],
reservoir_weight[146][193],
reservoir_weight[146][194],
reservoir_weight[146][195],
reservoir_weight[146][196],
reservoir_weight[146][197],
reservoir_weight[146][198],
reservoir_weight[146][199]
},
{reservoir_weight[147][0],
reservoir_weight[147][1],
reservoir_weight[147][2],
reservoir_weight[147][3],
reservoir_weight[147][4],
reservoir_weight[147][5],
reservoir_weight[147][6],
reservoir_weight[147][7],
reservoir_weight[147][8],
reservoir_weight[147][9],
reservoir_weight[147][10],
reservoir_weight[147][11],
reservoir_weight[147][12],
reservoir_weight[147][13],
reservoir_weight[147][14],
reservoir_weight[147][15],
reservoir_weight[147][16],
reservoir_weight[147][17],
reservoir_weight[147][18],
reservoir_weight[147][19],
reservoir_weight[147][20],
reservoir_weight[147][21],
reservoir_weight[147][22],
reservoir_weight[147][23],
reservoir_weight[147][24],
reservoir_weight[147][25],
reservoir_weight[147][26],
reservoir_weight[147][27],
reservoir_weight[147][28],
reservoir_weight[147][29],
reservoir_weight[147][30],
reservoir_weight[147][31],
reservoir_weight[147][32],
reservoir_weight[147][33],
reservoir_weight[147][34],
reservoir_weight[147][35],
reservoir_weight[147][36],
reservoir_weight[147][37],
reservoir_weight[147][38],
reservoir_weight[147][39],
reservoir_weight[147][40],
reservoir_weight[147][41],
reservoir_weight[147][42],
reservoir_weight[147][43],
reservoir_weight[147][44],
reservoir_weight[147][45],
reservoir_weight[147][46],
reservoir_weight[147][47],
reservoir_weight[147][48],
reservoir_weight[147][49],
reservoir_weight[147][50],
reservoir_weight[147][51],
reservoir_weight[147][52],
reservoir_weight[147][53],
reservoir_weight[147][54],
reservoir_weight[147][55],
reservoir_weight[147][56],
reservoir_weight[147][57],
reservoir_weight[147][58],
reservoir_weight[147][59],
reservoir_weight[147][60],
reservoir_weight[147][61],
reservoir_weight[147][62],
reservoir_weight[147][63],
reservoir_weight[147][64],
reservoir_weight[147][65],
reservoir_weight[147][66],
reservoir_weight[147][67],
reservoir_weight[147][68],
reservoir_weight[147][69],
reservoir_weight[147][70],
reservoir_weight[147][71],
reservoir_weight[147][72],
reservoir_weight[147][73],
reservoir_weight[147][74],
reservoir_weight[147][75],
reservoir_weight[147][76],
reservoir_weight[147][77],
reservoir_weight[147][78],
reservoir_weight[147][79],
reservoir_weight[147][80],
reservoir_weight[147][81],
reservoir_weight[147][82],
reservoir_weight[147][83],
reservoir_weight[147][84],
reservoir_weight[147][85],
reservoir_weight[147][86],
reservoir_weight[147][87],
reservoir_weight[147][88],
reservoir_weight[147][89],
reservoir_weight[147][90],
reservoir_weight[147][91],
reservoir_weight[147][92],
reservoir_weight[147][93],
reservoir_weight[147][94],
reservoir_weight[147][95],
reservoir_weight[147][96],
reservoir_weight[147][97],
reservoir_weight[147][98],
reservoir_weight[147][99],
reservoir_weight[147][100],
reservoir_weight[147][101],
reservoir_weight[147][102],
reservoir_weight[147][103],
reservoir_weight[147][104],
reservoir_weight[147][105],
reservoir_weight[147][106],
reservoir_weight[147][107],
reservoir_weight[147][108],
reservoir_weight[147][109],
reservoir_weight[147][110],
reservoir_weight[147][111],
reservoir_weight[147][112],
reservoir_weight[147][113],
reservoir_weight[147][114],
reservoir_weight[147][115],
reservoir_weight[147][116],
reservoir_weight[147][117],
reservoir_weight[147][118],
reservoir_weight[147][119],
reservoir_weight[147][120],
reservoir_weight[147][121],
reservoir_weight[147][122],
reservoir_weight[147][123],
reservoir_weight[147][124],
reservoir_weight[147][125],
reservoir_weight[147][126],
reservoir_weight[147][127],
reservoir_weight[147][128],
reservoir_weight[147][129],
reservoir_weight[147][130],
reservoir_weight[147][131],
reservoir_weight[147][132],
reservoir_weight[147][133],
reservoir_weight[147][134],
reservoir_weight[147][135],
reservoir_weight[147][136],
reservoir_weight[147][137],
reservoir_weight[147][138],
reservoir_weight[147][139],
reservoir_weight[147][140],
reservoir_weight[147][141],
reservoir_weight[147][142],
reservoir_weight[147][143],
reservoir_weight[147][144],
reservoir_weight[147][145],
reservoir_weight[147][146],
reservoir_weight[147][147],
reservoir_weight[147][148],
reservoir_weight[147][149],
reservoir_weight[147][150],
reservoir_weight[147][151],
reservoir_weight[147][152],
reservoir_weight[147][153],
reservoir_weight[147][154],
reservoir_weight[147][155],
reservoir_weight[147][156],
reservoir_weight[147][157],
reservoir_weight[147][158],
reservoir_weight[147][159],
reservoir_weight[147][160],
reservoir_weight[147][161],
reservoir_weight[147][162],
reservoir_weight[147][163],
reservoir_weight[147][164],
reservoir_weight[147][165],
reservoir_weight[147][166],
reservoir_weight[147][167],
reservoir_weight[147][168],
reservoir_weight[147][169],
reservoir_weight[147][170],
reservoir_weight[147][171],
reservoir_weight[147][172],
reservoir_weight[147][173],
reservoir_weight[147][174],
reservoir_weight[147][175],
reservoir_weight[147][176],
reservoir_weight[147][177],
reservoir_weight[147][178],
reservoir_weight[147][179],
reservoir_weight[147][180],
reservoir_weight[147][181],
reservoir_weight[147][182],
reservoir_weight[147][183],
reservoir_weight[147][184],
reservoir_weight[147][185],
reservoir_weight[147][186],
reservoir_weight[147][187],
reservoir_weight[147][188],
reservoir_weight[147][189],
reservoir_weight[147][190],
reservoir_weight[147][191],
reservoir_weight[147][192],
reservoir_weight[147][193],
reservoir_weight[147][194],
reservoir_weight[147][195],
reservoir_weight[147][196],
reservoir_weight[147][197],
reservoir_weight[147][198],
reservoir_weight[147][199]
},
{reservoir_weight[148][0],
reservoir_weight[148][1],
reservoir_weight[148][2],
reservoir_weight[148][3],
reservoir_weight[148][4],
reservoir_weight[148][5],
reservoir_weight[148][6],
reservoir_weight[148][7],
reservoir_weight[148][8],
reservoir_weight[148][9],
reservoir_weight[148][10],
reservoir_weight[148][11],
reservoir_weight[148][12],
reservoir_weight[148][13],
reservoir_weight[148][14],
reservoir_weight[148][15],
reservoir_weight[148][16],
reservoir_weight[148][17],
reservoir_weight[148][18],
reservoir_weight[148][19],
reservoir_weight[148][20],
reservoir_weight[148][21],
reservoir_weight[148][22],
reservoir_weight[148][23],
reservoir_weight[148][24],
reservoir_weight[148][25],
reservoir_weight[148][26],
reservoir_weight[148][27],
reservoir_weight[148][28],
reservoir_weight[148][29],
reservoir_weight[148][30],
reservoir_weight[148][31],
reservoir_weight[148][32],
reservoir_weight[148][33],
reservoir_weight[148][34],
reservoir_weight[148][35],
reservoir_weight[148][36],
reservoir_weight[148][37],
reservoir_weight[148][38],
reservoir_weight[148][39],
reservoir_weight[148][40],
reservoir_weight[148][41],
reservoir_weight[148][42],
reservoir_weight[148][43],
reservoir_weight[148][44],
reservoir_weight[148][45],
reservoir_weight[148][46],
reservoir_weight[148][47],
reservoir_weight[148][48],
reservoir_weight[148][49],
reservoir_weight[148][50],
reservoir_weight[148][51],
reservoir_weight[148][52],
reservoir_weight[148][53],
reservoir_weight[148][54],
reservoir_weight[148][55],
reservoir_weight[148][56],
reservoir_weight[148][57],
reservoir_weight[148][58],
reservoir_weight[148][59],
reservoir_weight[148][60],
reservoir_weight[148][61],
reservoir_weight[148][62],
reservoir_weight[148][63],
reservoir_weight[148][64],
reservoir_weight[148][65],
reservoir_weight[148][66],
reservoir_weight[148][67],
reservoir_weight[148][68],
reservoir_weight[148][69],
reservoir_weight[148][70],
reservoir_weight[148][71],
reservoir_weight[148][72],
reservoir_weight[148][73],
reservoir_weight[148][74],
reservoir_weight[148][75],
reservoir_weight[148][76],
reservoir_weight[148][77],
reservoir_weight[148][78],
reservoir_weight[148][79],
reservoir_weight[148][80],
reservoir_weight[148][81],
reservoir_weight[148][82],
reservoir_weight[148][83],
reservoir_weight[148][84],
reservoir_weight[148][85],
reservoir_weight[148][86],
reservoir_weight[148][87],
reservoir_weight[148][88],
reservoir_weight[148][89],
reservoir_weight[148][90],
reservoir_weight[148][91],
reservoir_weight[148][92],
reservoir_weight[148][93],
reservoir_weight[148][94],
reservoir_weight[148][95],
reservoir_weight[148][96],
reservoir_weight[148][97],
reservoir_weight[148][98],
reservoir_weight[148][99],
reservoir_weight[148][100],
reservoir_weight[148][101],
reservoir_weight[148][102],
reservoir_weight[148][103],
reservoir_weight[148][104],
reservoir_weight[148][105],
reservoir_weight[148][106],
reservoir_weight[148][107],
reservoir_weight[148][108],
reservoir_weight[148][109],
reservoir_weight[148][110],
reservoir_weight[148][111],
reservoir_weight[148][112],
reservoir_weight[148][113],
reservoir_weight[148][114],
reservoir_weight[148][115],
reservoir_weight[148][116],
reservoir_weight[148][117],
reservoir_weight[148][118],
reservoir_weight[148][119],
reservoir_weight[148][120],
reservoir_weight[148][121],
reservoir_weight[148][122],
reservoir_weight[148][123],
reservoir_weight[148][124],
reservoir_weight[148][125],
reservoir_weight[148][126],
reservoir_weight[148][127],
reservoir_weight[148][128],
reservoir_weight[148][129],
reservoir_weight[148][130],
reservoir_weight[148][131],
reservoir_weight[148][132],
reservoir_weight[148][133],
reservoir_weight[148][134],
reservoir_weight[148][135],
reservoir_weight[148][136],
reservoir_weight[148][137],
reservoir_weight[148][138],
reservoir_weight[148][139],
reservoir_weight[148][140],
reservoir_weight[148][141],
reservoir_weight[148][142],
reservoir_weight[148][143],
reservoir_weight[148][144],
reservoir_weight[148][145],
reservoir_weight[148][146],
reservoir_weight[148][147],
reservoir_weight[148][148],
reservoir_weight[148][149],
reservoir_weight[148][150],
reservoir_weight[148][151],
reservoir_weight[148][152],
reservoir_weight[148][153],
reservoir_weight[148][154],
reservoir_weight[148][155],
reservoir_weight[148][156],
reservoir_weight[148][157],
reservoir_weight[148][158],
reservoir_weight[148][159],
reservoir_weight[148][160],
reservoir_weight[148][161],
reservoir_weight[148][162],
reservoir_weight[148][163],
reservoir_weight[148][164],
reservoir_weight[148][165],
reservoir_weight[148][166],
reservoir_weight[148][167],
reservoir_weight[148][168],
reservoir_weight[148][169],
reservoir_weight[148][170],
reservoir_weight[148][171],
reservoir_weight[148][172],
reservoir_weight[148][173],
reservoir_weight[148][174],
reservoir_weight[148][175],
reservoir_weight[148][176],
reservoir_weight[148][177],
reservoir_weight[148][178],
reservoir_weight[148][179],
reservoir_weight[148][180],
reservoir_weight[148][181],
reservoir_weight[148][182],
reservoir_weight[148][183],
reservoir_weight[148][184],
reservoir_weight[148][185],
reservoir_weight[148][186],
reservoir_weight[148][187],
reservoir_weight[148][188],
reservoir_weight[148][189],
reservoir_weight[148][190],
reservoir_weight[148][191],
reservoir_weight[148][192],
reservoir_weight[148][193],
reservoir_weight[148][194],
reservoir_weight[148][195],
reservoir_weight[148][196],
reservoir_weight[148][197],
reservoir_weight[148][198],
reservoir_weight[148][199]
},
{reservoir_weight[149][0],
reservoir_weight[149][1],
reservoir_weight[149][2],
reservoir_weight[149][3],
reservoir_weight[149][4],
reservoir_weight[149][5],
reservoir_weight[149][6],
reservoir_weight[149][7],
reservoir_weight[149][8],
reservoir_weight[149][9],
reservoir_weight[149][10],
reservoir_weight[149][11],
reservoir_weight[149][12],
reservoir_weight[149][13],
reservoir_weight[149][14],
reservoir_weight[149][15],
reservoir_weight[149][16],
reservoir_weight[149][17],
reservoir_weight[149][18],
reservoir_weight[149][19],
reservoir_weight[149][20],
reservoir_weight[149][21],
reservoir_weight[149][22],
reservoir_weight[149][23],
reservoir_weight[149][24],
reservoir_weight[149][25],
reservoir_weight[149][26],
reservoir_weight[149][27],
reservoir_weight[149][28],
reservoir_weight[149][29],
reservoir_weight[149][30],
reservoir_weight[149][31],
reservoir_weight[149][32],
reservoir_weight[149][33],
reservoir_weight[149][34],
reservoir_weight[149][35],
reservoir_weight[149][36],
reservoir_weight[149][37],
reservoir_weight[149][38],
reservoir_weight[149][39],
reservoir_weight[149][40],
reservoir_weight[149][41],
reservoir_weight[149][42],
reservoir_weight[149][43],
reservoir_weight[149][44],
reservoir_weight[149][45],
reservoir_weight[149][46],
reservoir_weight[149][47],
reservoir_weight[149][48],
reservoir_weight[149][49],
reservoir_weight[149][50],
reservoir_weight[149][51],
reservoir_weight[149][52],
reservoir_weight[149][53],
reservoir_weight[149][54],
reservoir_weight[149][55],
reservoir_weight[149][56],
reservoir_weight[149][57],
reservoir_weight[149][58],
reservoir_weight[149][59],
reservoir_weight[149][60],
reservoir_weight[149][61],
reservoir_weight[149][62],
reservoir_weight[149][63],
reservoir_weight[149][64],
reservoir_weight[149][65],
reservoir_weight[149][66],
reservoir_weight[149][67],
reservoir_weight[149][68],
reservoir_weight[149][69],
reservoir_weight[149][70],
reservoir_weight[149][71],
reservoir_weight[149][72],
reservoir_weight[149][73],
reservoir_weight[149][74],
reservoir_weight[149][75],
reservoir_weight[149][76],
reservoir_weight[149][77],
reservoir_weight[149][78],
reservoir_weight[149][79],
reservoir_weight[149][80],
reservoir_weight[149][81],
reservoir_weight[149][82],
reservoir_weight[149][83],
reservoir_weight[149][84],
reservoir_weight[149][85],
reservoir_weight[149][86],
reservoir_weight[149][87],
reservoir_weight[149][88],
reservoir_weight[149][89],
reservoir_weight[149][90],
reservoir_weight[149][91],
reservoir_weight[149][92],
reservoir_weight[149][93],
reservoir_weight[149][94],
reservoir_weight[149][95],
reservoir_weight[149][96],
reservoir_weight[149][97],
reservoir_weight[149][98],
reservoir_weight[149][99],
reservoir_weight[149][100],
reservoir_weight[149][101],
reservoir_weight[149][102],
reservoir_weight[149][103],
reservoir_weight[149][104],
reservoir_weight[149][105],
reservoir_weight[149][106],
reservoir_weight[149][107],
reservoir_weight[149][108],
reservoir_weight[149][109],
reservoir_weight[149][110],
reservoir_weight[149][111],
reservoir_weight[149][112],
reservoir_weight[149][113],
reservoir_weight[149][114],
reservoir_weight[149][115],
reservoir_weight[149][116],
reservoir_weight[149][117],
reservoir_weight[149][118],
reservoir_weight[149][119],
reservoir_weight[149][120],
reservoir_weight[149][121],
reservoir_weight[149][122],
reservoir_weight[149][123],
reservoir_weight[149][124],
reservoir_weight[149][125],
reservoir_weight[149][126],
reservoir_weight[149][127],
reservoir_weight[149][128],
reservoir_weight[149][129],
reservoir_weight[149][130],
reservoir_weight[149][131],
reservoir_weight[149][132],
reservoir_weight[149][133],
reservoir_weight[149][134],
reservoir_weight[149][135],
reservoir_weight[149][136],
reservoir_weight[149][137],
reservoir_weight[149][138],
reservoir_weight[149][139],
reservoir_weight[149][140],
reservoir_weight[149][141],
reservoir_weight[149][142],
reservoir_weight[149][143],
reservoir_weight[149][144],
reservoir_weight[149][145],
reservoir_weight[149][146],
reservoir_weight[149][147],
reservoir_weight[149][148],
reservoir_weight[149][149],
reservoir_weight[149][150],
reservoir_weight[149][151],
reservoir_weight[149][152],
reservoir_weight[149][153],
reservoir_weight[149][154],
reservoir_weight[149][155],
reservoir_weight[149][156],
reservoir_weight[149][157],
reservoir_weight[149][158],
reservoir_weight[149][159],
reservoir_weight[149][160],
reservoir_weight[149][161],
reservoir_weight[149][162],
reservoir_weight[149][163],
reservoir_weight[149][164],
reservoir_weight[149][165],
reservoir_weight[149][166],
reservoir_weight[149][167],
reservoir_weight[149][168],
reservoir_weight[149][169],
reservoir_weight[149][170],
reservoir_weight[149][171],
reservoir_weight[149][172],
reservoir_weight[149][173],
reservoir_weight[149][174],
reservoir_weight[149][175],
reservoir_weight[149][176],
reservoir_weight[149][177],
reservoir_weight[149][178],
reservoir_weight[149][179],
reservoir_weight[149][180],
reservoir_weight[149][181],
reservoir_weight[149][182],
reservoir_weight[149][183],
reservoir_weight[149][184],
reservoir_weight[149][185],
reservoir_weight[149][186],
reservoir_weight[149][187],
reservoir_weight[149][188],
reservoir_weight[149][189],
reservoir_weight[149][190],
reservoir_weight[149][191],
reservoir_weight[149][192],
reservoir_weight[149][193],
reservoir_weight[149][194],
reservoir_weight[149][195],
reservoir_weight[149][196],
reservoir_weight[149][197],
reservoir_weight[149][198],
reservoir_weight[149][199]
},
{reservoir_weight[150][0],
reservoir_weight[150][1],
reservoir_weight[150][2],
reservoir_weight[150][3],
reservoir_weight[150][4],
reservoir_weight[150][5],
reservoir_weight[150][6],
reservoir_weight[150][7],
reservoir_weight[150][8],
reservoir_weight[150][9],
reservoir_weight[150][10],
reservoir_weight[150][11],
reservoir_weight[150][12],
reservoir_weight[150][13],
reservoir_weight[150][14],
reservoir_weight[150][15],
reservoir_weight[150][16],
reservoir_weight[150][17],
reservoir_weight[150][18],
reservoir_weight[150][19],
reservoir_weight[150][20],
reservoir_weight[150][21],
reservoir_weight[150][22],
reservoir_weight[150][23],
reservoir_weight[150][24],
reservoir_weight[150][25],
reservoir_weight[150][26],
reservoir_weight[150][27],
reservoir_weight[150][28],
reservoir_weight[150][29],
reservoir_weight[150][30],
reservoir_weight[150][31],
reservoir_weight[150][32],
reservoir_weight[150][33],
reservoir_weight[150][34],
reservoir_weight[150][35],
reservoir_weight[150][36],
reservoir_weight[150][37],
reservoir_weight[150][38],
reservoir_weight[150][39],
reservoir_weight[150][40],
reservoir_weight[150][41],
reservoir_weight[150][42],
reservoir_weight[150][43],
reservoir_weight[150][44],
reservoir_weight[150][45],
reservoir_weight[150][46],
reservoir_weight[150][47],
reservoir_weight[150][48],
reservoir_weight[150][49],
reservoir_weight[150][50],
reservoir_weight[150][51],
reservoir_weight[150][52],
reservoir_weight[150][53],
reservoir_weight[150][54],
reservoir_weight[150][55],
reservoir_weight[150][56],
reservoir_weight[150][57],
reservoir_weight[150][58],
reservoir_weight[150][59],
reservoir_weight[150][60],
reservoir_weight[150][61],
reservoir_weight[150][62],
reservoir_weight[150][63],
reservoir_weight[150][64],
reservoir_weight[150][65],
reservoir_weight[150][66],
reservoir_weight[150][67],
reservoir_weight[150][68],
reservoir_weight[150][69],
reservoir_weight[150][70],
reservoir_weight[150][71],
reservoir_weight[150][72],
reservoir_weight[150][73],
reservoir_weight[150][74],
reservoir_weight[150][75],
reservoir_weight[150][76],
reservoir_weight[150][77],
reservoir_weight[150][78],
reservoir_weight[150][79],
reservoir_weight[150][80],
reservoir_weight[150][81],
reservoir_weight[150][82],
reservoir_weight[150][83],
reservoir_weight[150][84],
reservoir_weight[150][85],
reservoir_weight[150][86],
reservoir_weight[150][87],
reservoir_weight[150][88],
reservoir_weight[150][89],
reservoir_weight[150][90],
reservoir_weight[150][91],
reservoir_weight[150][92],
reservoir_weight[150][93],
reservoir_weight[150][94],
reservoir_weight[150][95],
reservoir_weight[150][96],
reservoir_weight[150][97],
reservoir_weight[150][98],
reservoir_weight[150][99],
reservoir_weight[150][100],
reservoir_weight[150][101],
reservoir_weight[150][102],
reservoir_weight[150][103],
reservoir_weight[150][104],
reservoir_weight[150][105],
reservoir_weight[150][106],
reservoir_weight[150][107],
reservoir_weight[150][108],
reservoir_weight[150][109],
reservoir_weight[150][110],
reservoir_weight[150][111],
reservoir_weight[150][112],
reservoir_weight[150][113],
reservoir_weight[150][114],
reservoir_weight[150][115],
reservoir_weight[150][116],
reservoir_weight[150][117],
reservoir_weight[150][118],
reservoir_weight[150][119],
reservoir_weight[150][120],
reservoir_weight[150][121],
reservoir_weight[150][122],
reservoir_weight[150][123],
reservoir_weight[150][124],
reservoir_weight[150][125],
reservoir_weight[150][126],
reservoir_weight[150][127],
reservoir_weight[150][128],
reservoir_weight[150][129],
reservoir_weight[150][130],
reservoir_weight[150][131],
reservoir_weight[150][132],
reservoir_weight[150][133],
reservoir_weight[150][134],
reservoir_weight[150][135],
reservoir_weight[150][136],
reservoir_weight[150][137],
reservoir_weight[150][138],
reservoir_weight[150][139],
reservoir_weight[150][140],
reservoir_weight[150][141],
reservoir_weight[150][142],
reservoir_weight[150][143],
reservoir_weight[150][144],
reservoir_weight[150][145],
reservoir_weight[150][146],
reservoir_weight[150][147],
reservoir_weight[150][148],
reservoir_weight[150][149],
reservoir_weight[150][150],
reservoir_weight[150][151],
reservoir_weight[150][152],
reservoir_weight[150][153],
reservoir_weight[150][154],
reservoir_weight[150][155],
reservoir_weight[150][156],
reservoir_weight[150][157],
reservoir_weight[150][158],
reservoir_weight[150][159],
reservoir_weight[150][160],
reservoir_weight[150][161],
reservoir_weight[150][162],
reservoir_weight[150][163],
reservoir_weight[150][164],
reservoir_weight[150][165],
reservoir_weight[150][166],
reservoir_weight[150][167],
reservoir_weight[150][168],
reservoir_weight[150][169],
reservoir_weight[150][170],
reservoir_weight[150][171],
reservoir_weight[150][172],
reservoir_weight[150][173],
reservoir_weight[150][174],
reservoir_weight[150][175],
reservoir_weight[150][176],
reservoir_weight[150][177],
reservoir_weight[150][178],
reservoir_weight[150][179],
reservoir_weight[150][180],
reservoir_weight[150][181],
reservoir_weight[150][182],
reservoir_weight[150][183],
reservoir_weight[150][184],
reservoir_weight[150][185],
reservoir_weight[150][186],
reservoir_weight[150][187],
reservoir_weight[150][188],
reservoir_weight[150][189],
reservoir_weight[150][190],
reservoir_weight[150][191],
reservoir_weight[150][192],
reservoir_weight[150][193],
reservoir_weight[150][194],
reservoir_weight[150][195],
reservoir_weight[150][196],
reservoir_weight[150][197],
reservoir_weight[150][198],
reservoir_weight[150][199]
},
{reservoir_weight[151][0],
reservoir_weight[151][1],
reservoir_weight[151][2],
reservoir_weight[151][3],
reservoir_weight[151][4],
reservoir_weight[151][5],
reservoir_weight[151][6],
reservoir_weight[151][7],
reservoir_weight[151][8],
reservoir_weight[151][9],
reservoir_weight[151][10],
reservoir_weight[151][11],
reservoir_weight[151][12],
reservoir_weight[151][13],
reservoir_weight[151][14],
reservoir_weight[151][15],
reservoir_weight[151][16],
reservoir_weight[151][17],
reservoir_weight[151][18],
reservoir_weight[151][19],
reservoir_weight[151][20],
reservoir_weight[151][21],
reservoir_weight[151][22],
reservoir_weight[151][23],
reservoir_weight[151][24],
reservoir_weight[151][25],
reservoir_weight[151][26],
reservoir_weight[151][27],
reservoir_weight[151][28],
reservoir_weight[151][29],
reservoir_weight[151][30],
reservoir_weight[151][31],
reservoir_weight[151][32],
reservoir_weight[151][33],
reservoir_weight[151][34],
reservoir_weight[151][35],
reservoir_weight[151][36],
reservoir_weight[151][37],
reservoir_weight[151][38],
reservoir_weight[151][39],
reservoir_weight[151][40],
reservoir_weight[151][41],
reservoir_weight[151][42],
reservoir_weight[151][43],
reservoir_weight[151][44],
reservoir_weight[151][45],
reservoir_weight[151][46],
reservoir_weight[151][47],
reservoir_weight[151][48],
reservoir_weight[151][49],
reservoir_weight[151][50],
reservoir_weight[151][51],
reservoir_weight[151][52],
reservoir_weight[151][53],
reservoir_weight[151][54],
reservoir_weight[151][55],
reservoir_weight[151][56],
reservoir_weight[151][57],
reservoir_weight[151][58],
reservoir_weight[151][59],
reservoir_weight[151][60],
reservoir_weight[151][61],
reservoir_weight[151][62],
reservoir_weight[151][63],
reservoir_weight[151][64],
reservoir_weight[151][65],
reservoir_weight[151][66],
reservoir_weight[151][67],
reservoir_weight[151][68],
reservoir_weight[151][69],
reservoir_weight[151][70],
reservoir_weight[151][71],
reservoir_weight[151][72],
reservoir_weight[151][73],
reservoir_weight[151][74],
reservoir_weight[151][75],
reservoir_weight[151][76],
reservoir_weight[151][77],
reservoir_weight[151][78],
reservoir_weight[151][79],
reservoir_weight[151][80],
reservoir_weight[151][81],
reservoir_weight[151][82],
reservoir_weight[151][83],
reservoir_weight[151][84],
reservoir_weight[151][85],
reservoir_weight[151][86],
reservoir_weight[151][87],
reservoir_weight[151][88],
reservoir_weight[151][89],
reservoir_weight[151][90],
reservoir_weight[151][91],
reservoir_weight[151][92],
reservoir_weight[151][93],
reservoir_weight[151][94],
reservoir_weight[151][95],
reservoir_weight[151][96],
reservoir_weight[151][97],
reservoir_weight[151][98],
reservoir_weight[151][99],
reservoir_weight[151][100],
reservoir_weight[151][101],
reservoir_weight[151][102],
reservoir_weight[151][103],
reservoir_weight[151][104],
reservoir_weight[151][105],
reservoir_weight[151][106],
reservoir_weight[151][107],
reservoir_weight[151][108],
reservoir_weight[151][109],
reservoir_weight[151][110],
reservoir_weight[151][111],
reservoir_weight[151][112],
reservoir_weight[151][113],
reservoir_weight[151][114],
reservoir_weight[151][115],
reservoir_weight[151][116],
reservoir_weight[151][117],
reservoir_weight[151][118],
reservoir_weight[151][119],
reservoir_weight[151][120],
reservoir_weight[151][121],
reservoir_weight[151][122],
reservoir_weight[151][123],
reservoir_weight[151][124],
reservoir_weight[151][125],
reservoir_weight[151][126],
reservoir_weight[151][127],
reservoir_weight[151][128],
reservoir_weight[151][129],
reservoir_weight[151][130],
reservoir_weight[151][131],
reservoir_weight[151][132],
reservoir_weight[151][133],
reservoir_weight[151][134],
reservoir_weight[151][135],
reservoir_weight[151][136],
reservoir_weight[151][137],
reservoir_weight[151][138],
reservoir_weight[151][139],
reservoir_weight[151][140],
reservoir_weight[151][141],
reservoir_weight[151][142],
reservoir_weight[151][143],
reservoir_weight[151][144],
reservoir_weight[151][145],
reservoir_weight[151][146],
reservoir_weight[151][147],
reservoir_weight[151][148],
reservoir_weight[151][149],
reservoir_weight[151][150],
reservoir_weight[151][151],
reservoir_weight[151][152],
reservoir_weight[151][153],
reservoir_weight[151][154],
reservoir_weight[151][155],
reservoir_weight[151][156],
reservoir_weight[151][157],
reservoir_weight[151][158],
reservoir_weight[151][159],
reservoir_weight[151][160],
reservoir_weight[151][161],
reservoir_weight[151][162],
reservoir_weight[151][163],
reservoir_weight[151][164],
reservoir_weight[151][165],
reservoir_weight[151][166],
reservoir_weight[151][167],
reservoir_weight[151][168],
reservoir_weight[151][169],
reservoir_weight[151][170],
reservoir_weight[151][171],
reservoir_weight[151][172],
reservoir_weight[151][173],
reservoir_weight[151][174],
reservoir_weight[151][175],
reservoir_weight[151][176],
reservoir_weight[151][177],
reservoir_weight[151][178],
reservoir_weight[151][179],
reservoir_weight[151][180],
reservoir_weight[151][181],
reservoir_weight[151][182],
reservoir_weight[151][183],
reservoir_weight[151][184],
reservoir_weight[151][185],
reservoir_weight[151][186],
reservoir_weight[151][187],
reservoir_weight[151][188],
reservoir_weight[151][189],
reservoir_weight[151][190],
reservoir_weight[151][191],
reservoir_weight[151][192],
reservoir_weight[151][193],
reservoir_weight[151][194],
reservoir_weight[151][195],
reservoir_weight[151][196],
reservoir_weight[151][197],
reservoir_weight[151][198],
reservoir_weight[151][199]
},
{reservoir_weight[152][0],
reservoir_weight[152][1],
reservoir_weight[152][2],
reservoir_weight[152][3],
reservoir_weight[152][4],
reservoir_weight[152][5],
reservoir_weight[152][6],
reservoir_weight[152][7],
reservoir_weight[152][8],
reservoir_weight[152][9],
reservoir_weight[152][10],
reservoir_weight[152][11],
reservoir_weight[152][12],
reservoir_weight[152][13],
reservoir_weight[152][14],
reservoir_weight[152][15],
reservoir_weight[152][16],
reservoir_weight[152][17],
reservoir_weight[152][18],
reservoir_weight[152][19],
reservoir_weight[152][20],
reservoir_weight[152][21],
reservoir_weight[152][22],
reservoir_weight[152][23],
reservoir_weight[152][24],
reservoir_weight[152][25],
reservoir_weight[152][26],
reservoir_weight[152][27],
reservoir_weight[152][28],
reservoir_weight[152][29],
reservoir_weight[152][30],
reservoir_weight[152][31],
reservoir_weight[152][32],
reservoir_weight[152][33],
reservoir_weight[152][34],
reservoir_weight[152][35],
reservoir_weight[152][36],
reservoir_weight[152][37],
reservoir_weight[152][38],
reservoir_weight[152][39],
reservoir_weight[152][40],
reservoir_weight[152][41],
reservoir_weight[152][42],
reservoir_weight[152][43],
reservoir_weight[152][44],
reservoir_weight[152][45],
reservoir_weight[152][46],
reservoir_weight[152][47],
reservoir_weight[152][48],
reservoir_weight[152][49],
reservoir_weight[152][50],
reservoir_weight[152][51],
reservoir_weight[152][52],
reservoir_weight[152][53],
reservoir_weight[152][54],
reservoir_weight[152][55],
reservoir_weight[152][56],
reservoir_weight[152][57],
reservoir_weight[152][58],
reservoir_weight[152][59],
reservoir_weight[152][60],
reservoir_weight[152][61],
reservoir_weight[152][62],
reservoir_weight[152][63],
reservoir_weight[152][64],
reservoir_weight[152][65],
reservoir_weight[152][66],
reservoir_weight[152][67],
reservoir_weight[152][68],
reservoir_weight[152][69],
reservoir_weight[152][70],
reservoir_weight[152][71],
reservoir_weight[152][72],
reservoir_weight[152][73],
reservoir_weight[152][74],
reservoir_weight[152][75],
reservoir_weight[152][76],
reservoir_weight[152][77],
reservoir_weight[152][78],
reservoir_weight[152][79],
reservoir_weight[152][80],
reservoir_weight[152][81],
reservoir_weight[152][82],
reservoir_weight[152][83],
reservoir_weight[152][84],
reservoir_weight[152][85],
reservoir_weight[152][86],
reservoir_weight[152][87],
reservoir_weight[152][88],
reservoir_weight[152][89],
reservoir_weight[152][90],
reservoir_weight[152][91],
reservoir_weight[152][92],
reservoir_weight[152][93],
reservoir_weight[152][94],
reservoir_weight[152][95],
reservoir_weight[152][96],
reservoir_weight[152][97],
reservoir_weight[152][98],
reservoir_weight[152][99],
reservoir_weight[152][100],
reservoir_weight[152][101],
reservoir_weight[152][102],
reservoir_weight[152][103],
reservoir_weight[152][104],
reservoir_weight[152][105],
reservoir_weight[152][106],
reservoir_weight[152][107],
reservoir_weight[152][108],
reservoir_weight[152][109],
reservoir_weight[152][110],
reservoir_weight[152][111],
reservoir_weight[152][112],
reservoir_weight[152][113],
reservoir_weight[152][114],
reservoir_weight[152][115],
reservoir_weight[152][116],
reservoir_weight[152][117],
reservoir_weight[152][118],
reservoir_weight[152][119],
reservoir_weight[152][120],
reservoir_weight[152][121],
reservoir_weight[152][122],
reservoir_weight[152][123],
reservoir_weight[152][124],
reservoir_weight[152][125],
reservoir_weight[152][126],
reservoir_weight[152][127],
reservoir_weight[152][128],
reservoir_weight[152][129],
reservoir_weight[152][130],
reservoir_weight[152][131],
reservoir_weight[152][132],
reservoir_weight[152][133],
reservoir_weight[152][134],
reservoir_weight[152][135],
reservoir_weight[152][136],
reservoir_weight[152][137],
reservoir_weight[152][138],
reservoir_weight[152][139],
reservoir_weight[152][140],
reservoir_weight[152][141],
reservoir_weight[152][142],
reservoir_weight[152][143],
reservoir_weight[152][144],
reservoir_weight[152][145],
reservoir_weight[152][146],
reservoir_weight[152][147],
reservoir_weight[152][148],
reservoir_weight[152][149],
reservoir_weight[152][150],
reservoir_weight[152][151],
reservoir_weight[152][152],
reservoir_weight[152][153],
reservoir_weight[152][154],
reservoir_weight[152][155],
reservoir_weight[152][156],
reservoir_weight[152][157],
reservoir_weight[152][158],
reservoir_weight[152][159],
reservoir_weight[152][160],
reservoir_weight[152][161],
reservoir_weight[152][162],
reservoir_weight[152][163],
reservoir_weight[152][164],
reservoir_weight[152][165],
reservoir_weight[152][166],
reservoir_weight[152][167],
reservoir_weight[152][168],
reservoir_weight[152][169],
reservoir_weight[152][170],
reservoir_weight[152][171],
reservoir_weight[152][172],
reservoir_weight[152][173],
reservoir_weight[152][174],
reservoir_weight[152][175],
reservoir_weight[152][176],
reservoir_weight[152][177],
reservoir_weight[152][178],
reservoir_weight[152][179],
reservoir_weight[152][180],
reservoir_weight[152][181],
reservoir_weight[152][182],
reservoir_weight[152][183],
reservoir_weight[152][184],
reservoir_weight[152][185],
reservoir_weight[152][186],
reservoir_weight[152][187],
reservoir_weight[152][188],
reservoir_weight[152][189],
reservoir_weight[152][190],
reservoir_weight[152][191],
reservoir_weight[152][192],
reservoir_weight[152][193],
reservoir_weight[152][194],
reservoir_weight[152][195],
reservoir_weight[152][196],
reservoir_weight[152][197],
reservoir_weight[152][198],
reservoir_weight[152][199]
},
{reservoir_weight[153][0],
reservoir_weight[153][1],
reservoir_weight[153][2],
reservoir_weight[153][3],
reservoir_weight[153][4],
reservoir_weight[153][5],
reservoir_weight[153][6],
reservoir_weight[153][7],
reservoir_weight[153][8],
reservoir_weight[153][9],
reservoir_weight[153][10],
reservoir_weight[153][11],
reservoir_weight[153][12],
reservoir_weight[153][13],
reservoir_weight[153][14],
reservoir_weight[153][15],
reservoir_weight[153][16],
reservoir_weight[153][17],
reservoir_weight[153][18],
reservoir_weight[153][19],
reservoir_weight[153][20],
reservoir_weight[153][21],
reservoir_weight[153][22],
reservoir_weight[153][23],
reservoir_weight[153][24],
reservoir_weight[153][25],
reservoir_weight[153][26],
reservoir_weight[153][27],
reservoir_weight[153][28],
reservoir_weight[153][29],
reservoir_weight[153][30],
reservoir_weight[153][31],
reservoir_weight[153][32],
reservoir_weight[153][33],
reservoir_weight[153][34],
reservoir_weight[153][35],
reservoir_weight[153][36],
reservoir_weight[153][37],
reservoir_weight[153][38],
reservoir_weight[153][39],
reservoir_weight[153][40],
reservoir_weight[153][41],
reservoir_weight[153][42],
reservoir_weight[153][43],
reservoir_weight[153][44],
reservoir_weight[153][45],
reservoir_weight[153][46],
reservoir_weight[153][47],
reservoir_weight[153][48],
reservoir_weight[153][49],
reservoir_weight[153][50],
reservoir_weight[153][51],
reservoir_weight[153][52],
reservoir_weight[153][53],
reservoir_weight[153][54],
reservoir_weight[153][55],
reservoir_weight[153][56],
reservoir_weight[153][57],
reservoir_weight[153][58],
reservoir_weight[153][59],
reservoir_weight[153][60],
reservoir_weight[153][61],
reservoir_weight[153][62],
reservoir_weight[153][63],
reservoir_weight[153][64],
reservoir_weight[153][65],
reservoir_weight[153][66],
reservoir_weight[153][67],
reservoir_weight[153][68],
reservoir_weight[153][69],
reservoir_weight[153][70],
reservoir_weight[153][71],
reservoir_weight[153][72],
reservoir_weight[153][73],
reservoir_weight[153][74],
reservoir_weight[153][75],
reservoir_weight[153][76],
reservoir_weight[153][77],
reservoir_weight[153][78],
reservoir_weight[153][79],
reservoir_weight[153][80],
reservoir_weight[153][81],
reservoir_weight[153][82],
reservoir_weight[153][83],
reservoir_weight[153][84],
reservoir_weight[153][85],
reservoir_weight[153][86],
reservoir_weight[153][87],
reservoir_weight[153][88],
reservoir_weight[153][89],
reservoir_weight[153][90],
reservoir_weight[153][91],
reservoir_weight[153][92],
reservoir_weight[153][93],
reservoir_weight[153][94],
reservoir_weight[153][95],
reservoir_weight[153][96],
reservoir_weight[153][97],
reservoir_weight[153][98],
reservoir_weight[153][99],
reservoir_weight[153][100],
reservoir_weight[153][101],
reservoir_weight[153][102],
reservoir_weight[153][103],
reservoir_weight[153][104],
reservoir_weight[153][105],
reservoir_weight[153][106],
reservoir_weight[153][107],
reservoir_weight[153][108],
reservoir_weight[153][109],
reservoir_weight[153][110],
reservoir_weight[153][111],
reservoir_weight[153][112],
reservoir_weight[153][113],
reservoir_weight[153][114],
reservoir_weight[153][115],
reservoir_weight[153][116],
reservoir_weight[153][117],
reservoir_weight[153][118],
reservoir_weight[153][119],
reservoir_weight[153][120],
reservoir_weight[153][121],
reservoir_weight[153][122],
reservoir_weight[153][123],
reservoir_weight[153][124],
reservoir_weight[153][125],
reservoir_weight[153][126],
reservoir_weight[153][127],
reservoir_weight[153][128],
reservoir_weight[153][129],
reservoir_weight[153][130],
reservoir_weight[153][131],
reservoir_weight[153][132],
reservoir_weight[153][133],
reservoir_weight[153][134],
reservoir_weight[153][135],
reservoir_weight[153][136],
reservoir_weight[153][137],
reservoir_weight[153][138],
reservoir_weight[153][139],
reservoir_weight[153][140],
reservoir_weight[153][141],
reservoir_weight[153][142],
reservoir_weight[153][143],
reservoir_weight[153][144],
reservoir_weight[153][145],
reservoir_weight[153][146],
reservoir_weight[153][147],
reservoir_weight[153][148],
reservoir_weight[153][149],
reservoir_weight[153][150],
reservoir_weight[153][151],
reservoir_weight[153][152],
reservoir_weight[153][153],
reservoir_weight[153][154],
reservoir_weight[153][155],
reservoir_weight[153][156],
reservoir_weight[153][157],
reservoir_weight[153][158],
reservoir_weight[153][159],
reservoir_weight[153][160],
reservoir_weight[153][161],
reservoir_weight[153][162],
reservoir_weight[153][163],
reservoir_weight[153][164],
reservoir_weight[153][165],
reservoir_weight[153][166],
reservoir_weight[153][167],
reservoir_weight[153][168],
reservoir_weight[153][169],
reservoir_weight[153][170],
reservoir_weight[153][171],
reservoir_weight[153][172],
reservoir_weight[153][173],
reservoir_weight[153][174],
reservoir_weight[153][175],
reservoir_weight[153][176],
reservoir_weight[153][177],
reservoir_weight[153][178],
reservoir_weight[153][179],
reservoir_weight[153][180],
reservoir_weight[153][181],
reservoir_weight[153][182],
reservoir_weight[153][183],
reservoir_weight[153][184],
reservoir_weight[153][185],
reservoir_weight[153][186],
reservoir_weight[153][187],
reservoir_weight[153][188],
reservoir_weight[153][189],
reservoir_weight[153][190],
reservoir_weight[153][191],
reservoir_weight[153][192],
reservoir_weight[153][193],
reservoir_weight[153][194],
reservoir_weight[153][195],
reservoir_weight[153][196],
reservoir_weight[153][197],
reservoir_weight[153][198],
reservoir_weight[153][199]
},
{reservoir_weight[154][0],
reservoir_weight[154][1],
reservoir_weight[154][2],
reservoir_weight[154][3],
reservoir_weight[154][4],
reservoir_weight[154][5],
reservoir_weight[154][6],
reservoir_weight[154][7],
reservoir_weight[154][8],
reservoir_weight[154][9],
reservoir_weight[154][10],
reservoir_weight[154][11],
reservoir_weight[154][12],
reservoir_weight[154][13],
reservoir_weight[154][14],
reservoir_weight[154][15],
reservoir_weight[154][16],
reservoir_weight[154][17],
reservoir_weight[154][18],
reservoir_weight[154][19],
reservoir_weight[154][20],
reservoir_weight[154][21],
reservoir_weight[154][22],
reservoir_weight[154][23],
reservoir_weight[154][24],
reservoir_weight[154][25],
reservoir_weight[154][26],
reservoir_weight[154][27],
reservoir_weight[154][28],
reservoir_weight[154][29],
reservoir_weight[154][30],
reservoir_weight[154][31],
reservoir_weight[154][32],
reservoir_weight[154][33],
reservoir_weight[154][34],
reservoir_weight[154][35],
reservoir_weight[154][36],
reservoir_weight[154][37],
reservoir_weight[154][38],
reservoir_weight[154][39],
reservoir_weight[154][40],
reservoir_weight[154][41],
reservoir_weight[154][42],
reservoir_weight[154][43],
reservoir_weight[154][44],
reservoir_weight[154][45],
reservoir_weight[154][46],
reservoir_weight[154][47],
reservoir_weight[154][48],
reservoir_weight[154][49],
reservoir_weight[154][50],
reservoir_weight[154][51],
reservoir_weight[154][52],
reservoir_weight[154][53],
reservoir_weight[154][54],
reservoir_weight[154][55],
reservoir_weight[154][56],
reservoir_weight[154][57],
reservoir_weight[154][58],
reservoir_weight[154][59],
reservoir_weight[154][60],
reservoir_weight[154][61],
reservoir_weight[154][62],
reservoir_weight[154][63],
reservoir_weight[154][64],
reservoir_weight[154][65],
reservoir_weight[154][66],
reservoir_weight[154][67],
reservoir_weight[154][68],
reservoir_weight[154][69],
reservoir_weight[154][70],
reservoir_weight[154][71],
reservoir_weight[154][72],
reservoir_weight[154][73],
reservoir_weight[154][74],
reservoir_weight[154][75],
reservoir_weight[154][76],
reservoir_weight[154][77],
reservoir_weight[154][78],
reservoir_weight[154][79],
reservoir_weight[154][80],
reservoir_weight[154][81],
reservoir_weight[154][82],
reservoir_weight[154][83],
reservoir_weight[154][84],
reservoir_weight[154][85],
reservoir_weight[154][86],
reservoir_weight[154][87],
reservoir_weight[154][88],
reservoir_weight[154][89],
reservoir_weight[154][90],
reservoir_weight[154][91],
reservoir_weight[154][92],
reservoir_weight[154][93],
reservoir_weight[154][94],
reservoir_weight[154][95],
reservoir_weight[154][96],
reservoir_weight[154][97],
reservoir_weight[154][98],
reservoir_weight[154][99],
reservoir_weight[154][100],
reservoir_weight[154][101],
reservoir_weight[154][102],
reservoir_weight[154][103],
reservoir_weight[154][104],
reservoir_weight[154][105],
reservoir_weight[154][106],
reservoir_weight[154][107],
reservoir_weight[154][108],
reservoir_weight[154][109],
reservoir_weight[154][110],
reservoir_weight[154][111],
reservoir_weight[154][112],
reservoir_weight[154][113],
reservoir_weight[154][114],
reservoir_weight[154][115],
reservoir_weight[154][116],
reservoir_weight[154][117],
reservoir_weight[154][118],
reservoir_weight[154][119],
reservoir_weight[154][120],
reservoir_weight[154][121],
reservoir_weight[154][122],
reservoir_weight[154][123],
reservoir_weight[154][124],
reservoir_weight[154][125],
reservoir_weight[154][126],
reservoir_weight[154][127],
reservoir_weight[154][128],
reservoir_weight[154][129],
reservoir_weight[154][130],
reservoir_weight[154][131],
reservoir_weight[154][132],
reservoir_weight[154][133],
reservoir_weight[154][134],
reservoir_weight[154][135],
reservoir_weight[154][136],
reservoir_weight[154][137],
reservoir_weight[154][138],
reservoir_weight[154][139],
reservoir_weight[154][140],
reservoir_weight[154][141],
reservoir_weight[154][142],
reservoir_weight[154][143],
reservoir_weight[154][144],
reservoir_weight[154][145],
reservoir_weight[154][146],
reservoir_weight[154][147],
reservoir_weight[154][148],
reservoir_weight[154][149],
reservoir_weight[154][150],
reservoir_weight[154][151],
reservoir_weight[154][152],
reservoir_weight[154][153],
reservoir_weight[154][154],
reservoir_weight[154][155],
reservoir_weight[154][156],
reservoir_weight[154][157],
reservoir_weight[154][158],
reservoir_weight[154][159],
reservoir_weight[154][160],
reservoir_weight[154][161],
reservoir_weight[154][162],
reservoir_weight[154][163],
reservoir_weight[154][164],
reservoir_weight[154][165],
reservoir_weight[154][166],
reservoir_weight[154][167],
reservoir_weight[154][168],
reservoir_weight[154][169],
reservoir_weight[154][170],
reservoir_weight[154][171],
reservoir_weight[154][172],
reservoir_weight[154][173],
reservoir_weight[154][174],
reservoir_weight[154][175],
reservoir_weight[154][176],
reservoir_weight[154][177],
reservoir_weight[154][178],
reservoir_weight[154][179],
reservoir_weight[154][180],
reservoir_weight[154][181],
reservoir_weight[154][182],
reservoir_weight[154][183],
reservoir_weight[154][184],
reservoir_weight[154][185],
reservoir_weight[154][186],
reservoir_weight[154][187],
reservoir_weight[154][188],
reservoir_weight[154][189],
reservoir_weight[154][190],
reservoir_weight[154][191],
reservoir_weight[154][192],
reservoir_weight[154][193],
reservoir_weight[154][194],
reservoir_weight[154][195],
reservoir_weight[154][196],
reservoir_weight[154][197],
reservoir_weight[154][198],
reservoir_weight[154][199]
},
{reservoir_weight[155][0],
reservoir_weight[155][1],
reservoir_weight[155][2],
reservoir_weight[155][3],
reservoir_weight[155][4],
reservoir_weight[155][5],
reservoir_weight[155][6],
reservoir_weight[155][7],
reservoir_weight[155][8],
reservoir_weight[155][9],
reservoir_weight[155][10],
reservoir_weight[155][11],
reservoir_weight[155][12],
reservoir_weight[155][13],
reservoir_weight[155][14],
reservoir_weight[155][15],
reservoir_weight[155][16],
reservoir_weight[155][17],
reservoir_weight[155][18],
reservoir_weight[155][19],
reservoir_weight[155][20],
reservoir_weight[155][21],
reservoir_weight[155][22],
reservoir_weight[155][23],
reservoir_weight[155][24],
reservoir_weight[155][25],
reservoir_weight[155][26],
reservoir_weight[155][27],
reservoir_weight[155][28],
reservoir_weight[155][29],
reservoir_weight[155][30],
reservoir_weight[155][31],
reservoir_weight[155][32],
reservoir_weight[155][33],
reservoir_weight[155][34],
reservoir_weight[155][35],
reservoir_weight[155][36],
reservoir_weight[155][37],
reservoir_weight[155][38],
reservoir_weight[155][39],
reservoir_weight[155][40],
reservoir_weight[155][41],
reservoir_weight[155][42],
reservoir_weight[155][43],
reservoir_weight[155][44],
reservoir_weight[155][45],
reservoir_weight[155][46],
reservoir_weight[155][47],
reservoir_weight[155][48],
reservoir_weight[155][49],
reservoir_weight[155][50],
reservoir_weight[155][51],
reservoir_weight[155][52],
reservoir_weight[155][53],
reservoir_weight[155][54],
reservoir_weight[155][55],
reservoir_weight[155][56],
reservoir_weight[155][57],
reservoir_weight[155][58],
reservoir_weight[155][59],
reservoir_weight[155][60],
reservoir_weight[155][61],
reservoir_weight[155][62],
reservoir_weight[155][63],
reservoir_weight[155][64],
reservoir_weight[155][65],
reservoir_weight[155][66],
reservoir_weight[155][67],
reservoir_weight[155][68],
reservoir_weight[155][69],
reservoir_weight[155][70],
reservoir_weight[155][71],
reservoir_weight[155][72],
reservoir_weight[155][73],
reservoir_weight[155][74],
reservoir_weight[155][75],
reservoir_weight[155][76],
reservoir_weight[155][77],
reservoir_weight[155][78],
reservoir_weight[155][79],
reservoir_weight[155][80],
reservoir_weight[155][81],
reservoir_weight[155][82],
reservoir_weight[155][83],
reservoir_weight[155][84],
reservoir_weight[155][85],
reservoir_weight[155][86],
reservoir_weight[155][87],
reservoir_weight[155][88],
reservoir_weight[155][89],
reservoir_weight[155][90],
reservoir_weight[155][91],
reservoir_weight[155][92],
reservoir_weight[155][93],
reservoir_weight[155][94],
reservoir_weight[155][95],
reservoir_weight[155][96],
reservoir_weight[155][97],
reservoir_weight[155][98],
reservoir_weight[155][99],
reservoir_weight[155][100],
reservoir_weight[155][101],
reservoir_weight[155][102],
reservoir_weight[155][103],
reservoir_weight[155][104],
reservoir_weight[155][105],
reservoir_weight[155][106],
reservoir_weight[155][107],
reservoir_weight[155][108],
reservoir_weight[155][109],
reservoir_weight[155][110],
reservoir_weight[155][111],
reservoir_weight[155][112],
reservoir_weight[155][113],
reservoir_weight[155][114],
reservoir_weight[155][115],
reservoir_weight[155][116],
reservoir_weight[155][117],
reservoir_weight[155][118],
reservoir_weight[155][119],
reservoir_weight[155][120],
reservoir_weight[155][121],
reservoir_weight[155][122],
reservoir_weight[155][123],
reservoir_weight[155][124],
reservoir_weight[155][125],
reservoir_weight[155][126],
reservoir_weight[155][127],
reservoir_weight[155][128],
reservoir_weight[155][129],
reservoir_weight[155][130],
reservoir_weight[155][131],
reservoir_weight[155][132],
reservoir_weight[155][133],
reservoir_weight[155][134],
reservoir_weight[155][135],
reservoir_weight[155][136],
reservoir_weight[155][137],
reservoir_weight[155][138],
reservoir_weight[155][139],
reservoir_weight[155][140],
reservoir_weight[155][141],
reservoir_weight[155][142],
reservoir_weight[155][143],
reservoir_weight[155][144],
reservoir_weight[155][145],
reservoir_weight[155][146],
reservoir_weight[155][147],
reservoir_weight[155][148],
reservoir_weight[155][149],
reservoir_weight[155][150],
reservoir_weight[155][151],
reservoir_weight[155][152],
reservoir_weight[155][153],
reservoir_weight[155][154],
reservoir_weight[155][155],
reservoir_weight[155][156],
reservoir_weight[155][157],
reservoir_weight[155][158],
reservoir_weight[155][159],
reservoir_weight[155][160],
reservoir_weight[155][161],
reservoir_weight[155][162],
reservoir_weight[155][163],
reservoir_weight[155][164],
reservoir_weight[155][165],
reservoir_weight[155][166],
reservoir_weight[155][167],
reservoir_weight[155][168],
reservoir_weight[155][169],
reservoir_weight[155][170],
reservoir_weight[155][171],
reservoir_weight[155][172],
reservoir_weight[155][173],
reservoir_weight[155][174],
reservoir_weight[155][175],
reservoir_weight[155][176],
reservoir_weight[155][177],
reservoir_weight[155][178],
reservoir_weight[155][179],
reservoir_weight[155][180],
reservoir_weight[155][181],
reservoir_weight[155][182],
reservoir_weight[155][183],
reservoir_weight[155][184],
reservoir_weight[155][185],
reservoir_weight[155][186],
reservoir_weight[155][187],
reservoir_weight[155][188],
reservoir_weight[155][189],
reservoir_weight[155][190],
reservoir_weight[155][191],
reservoir_weight[155][192],
reservoir_weight[155][193],
reservoir_weight[155][194],
reservoir_weight[155][195],
reservoir_weight[155][196],
reservoir_weight[155][197],
reservoir_weight[155][198],
reservoir_weight[155][199]
},
{reservoir_weight[156][0],
reservoir_weight[156][1],
reservoir_weight[156][2],
reservoir_weight[156][3],
reservoir_weight[156][4],
reservoir_weight[156][5],
reservoir_weight[156][6],
reservoir_weight[156][7],
reservoir_weight[156][8],
reservoir_weight[156][9],
reservoir_weight[156][10],
reservoir_weight[156][11],
reservoir_weight[156][12],
reservoir_weight[156][13],
reservoir_weight[156][14],
reservoir_weight[156][15],
reservoir_weight[156][16],
reservoir_weight[156][17],
reservoir_weight[156][18],
reservoir_weight[156][19],
reservoir_weight[156][20],
reservoir_weight[156][21],
reservoir_weight[156][22],
reservoir_weight[156][23],
reservoir_weight[156][24],
reservoir_weight[156][25],
reservoir_weight[156][26],
reservoir_weight[156][27],
reservoir_weight[156][28],
reservoir_weight[156][29],
reservoir_weight[156][30],
reservoir_weight[156][31],
reservoir_weight[156][32],
reservoir_weight[156][33],
reservoir_weight[156][34],
reservoir_weight[156][35],
reservoir_weight[156][36],
reservoir_weight[156][37],
reservoir_weight[156][38],
reservoir_weight[156][39],
reservoir_weight[156][40],
reservoir_weight[156][41],
reservoir_weight[156][42],
reservoir_weight[156][43],
reservoir_weight[156][44],
reservoir_weight[156][45],
reservoir_weight[156][46],
reservoir_weight[156][47],
reservoir_weight[156][48],
reservoir_weight[156][49],
reservoir_weight[156][50],
reservoir_weight[156][51],
reservoir_weight[156][52],
reservoir_weight[156][53],
reservoir_weight[156][54],
reservoir_weight[156][55],
reservoir_weight[156][56],
reservoir_weight[156][57],
reservoir_weight[156][58],
reservoir_weight[156][59],
reservoir_weight[156][60],
reservoir_weight[156][61],
reservoir_weight[156][62],
reservoir_weight[156][63],
reservoir_weight[156][64],
reservoir_weight[156][65],
reservoir_weight[156][66],
reservoir_weight[156][67],
reservoir_weight[156][68],
reservoir_weight[156][69],
reservoir_weight[156][70],
reservoir_weight[156][71],
reservoir_weight[156][72],
reservoir_weight[156][73],
reservoir_weight[156][74],
reservoir_weight[156][75],
reservoir_weight[156][76],
reservoir_weight[156][77],
reservoir_weight[156][78],
reservoir_weight[156][79],
reservoir_weight[156][80],
reservoir_weight[156][81],
reservoir_weight[156][82],
reservoir_weight[156][83],
reservoir_weight[156][84],
reservoir_weight[156][85],
reservoir_weight[156][86],
reservoir_weight[156][87],
reservoir_weight[156][88],
reservoir_weight[156][89],
reservoir_weight[156][90],
reservoir_weight[156][91],
reservoir_weight[156][92],
reservoir_weight[156][93],
reservoir_weight[156][94],
reservoir_weight[156][95],
reservoir_weight[156][96],
reservoir_weight[156][97],
reservoir_weight[156][98],
reservoir_weight[156][99],
reservoir_weight[156][100],
reservoir_weight[156][101],
reservoir_weight[156][102],
reservoir_weight[156][103],
reservoir_weight[156][104],
reservoir_weight[156][105],
reservoir_weight[156][106],
reservoir_weight[156][107],
reservoir_weight[156][108],
reservoir_weight[156][109],
reservoir_weight[156][110],
reservoir_weight[156][111],
reservoir_weight[156][112],
reservoir_weight[156][113],
reservoir_weight[156][114],
reservoir_weight[156][115],
reservoir_weight[156][116],
reservoir_weight[156][117],
reservoir_weight[156][118],
reservoir_weight[156][119],
reservoir_weight[156][120],
reservoir_weight[156][121],
reservoir_weight[156][122],
reservoir_weight[156][123],
reservoir_weight[156][124],
reservoir_weight[156][125],
reservoir_weight[156][126],
reservoir_weight[156][127],
reservoir_weight[156][128],
reservoir_weight[156][129],
reservoir_weight[156][130],
reservoir_weight[156][131],
reservoir_weight[156][132],
reservoir_weight[156][133],
reservoir_weight[156][134],
reservoir_weight[156][135],
reservoir_weight[156][136],
reservoir_weight[156][137],
reservoir_weight[156][138],
reservoir_weight[156][139],
reservoir_weight[156][140],
reservoir_weight[156][141],
reservoir_weight[156][142],
reservoir_weight[156][143],
reservoir_weight[156][144],
reservoir_weight[156][145],
reservoir_weight[156][146],
reservoir_weight[156][147],
reservoir_weight[156][148],
reservoir_weight[156][149],
reservoir_weight[156][150],
reservoir_weight[156][151],
reservoir_weight[156][152],
reservoir_weight[156][153],
reservoir_weight[156][154],
reservoir_weight[156][155],
reservoir_weight[156][156],
reservoir_weight[156][157],
reservoir_weight[156][158],
reservoir_weight[156][159],
reservoir_weight[156][160],
reservoir_weight[156][161],
reservoir_weight[156][162],
reservoir_weight[156][163],
reservoir_weight[156][164],
reservoir_weight[156][165],
reservoir_weight[156][166],
reservoir_weight[156][167],
reservoir_weight[156][168],
reservoir_weight[156][169],
reservoir_weight[156][170],
reservoir_weight[156][171],
reservoir_weight[156][172],
reservoir_weight[156][173],
reservoir_weight[156][174],
reservoir_weight[156][175],
reservoir_weight[156][176],
reservoir_weight[156][177],
reservoir_weight[156][178],
reservoir_weight[156][179],
reservoir_weight[156][180],
reservoir_weight[156][181],
reservoir_weight[156][182],
reservoir_weight[156][183],
reservoir_weight[156][184],
reservoir_weight[156][185],
reservoir_weight[156][186],
reservoir_weight[156][187],
reservoir_weight[156][188],
reservoir_weight[156][189],
reservoir_weight[156][190],
reservoir_weight[156][191],
reservoir_weight[156][192],
reservoir_weight[156][193],
reservoir_weight[156][194],
reservoir_weight[156][195],
reservoir_weight[156][196],
reservoir_weight[156][197],
reservoir_weight[156][198],
reservoir_weight[156][199]
},
{reservoir_weight[157][0],
reservoir_weight[157][1],
reservoir_weight[157][2],
reservoir_weight[157][3],
reservoir_weight[157][4],
reservoir_weight[157][5],
reservoir_weight[157][6],
reservoir_weight[157][7],
reservoir_weight[157][8],
reservoir_weight[157][9],
reservoir_weight[157][10],
reservoir_weight[157][11],
reservoir_weight[157][12],
reservoir_weight[157][13],
reservoir_weight[157][14],
reservoir_weight[157][15],
reservoir_weight[157][16],
reservoir_weight[157][17],
reservoir_weight[157][18],
reservoir_weight[157][19],
reservoir_weight[157][20],
reservoir_weight[157][21],
reservoir_weight[157][22],
reservoir_weight[157][23],
reservoir_weight[157][24],
reservoir_weight[157][25],
reservoir_weight[157][26],
reservoir_weight[157][27],
reservoir_weight[157][28],
reservoir_weight[157][29],
reservoir_weight[157][30],
reservoir_weight[157][31],
reservoir_weight[157][32],
reservoir_weight[157][33],
reservoir_weight[157][34],
reservoir_weight[157][35],
reservoir_weight[157][36],
reservoir_weight[157][37],
reservoir_weight[157][38],
reservoir_weight[157][39],
reservoir_weight[157][40],
reservoir_weight[157][41],
reservoir_weight[157][42],
reservoir_weight[157][43],
reservoir_weight[157][44],
reservoir_weight[157][45],
reservoir_weight[157][46],
reservoir_weight[157][47],
reservoir_weight[157][48],
reservoir_weight[157][49],
reservoir_weight[157][50],
reservoir_weight[157][51],
reservoir_weight[157][52],
reservoir_weight[157][53],
reservoir_weight[157][54],
reservoir_weight[157][55],
reservoir_weight[157][56],
reservoir_weight[157][57],
reservoir_weight[157][58],
reservoir_weight[157][59],
reservoir_weight[157][60],
reservoir_weight[157][61],
reservoir_weight[157][62],
reservoir_weight[157][63],
reservoir_weight[157][64],
reservoir_weight[157][65],
reservoir_weight[157][66],
reservoir_weight[157][67],
reservoir_weight[157][68],
reservoir_weight[157][69],
reservoir_weight[157][70],
reservoir_weight[157][71],
reservoir_weight[157][72],
reservoir_weight[157][73],
reservoir_weight[157][74],
reservoir_weight[157][75],
reservoir_weight[157][76],
reservoir_weight[157][77],
reservoir_weight[157][78],
reservoir_weight[157][79],
reservoir_weight[157][80],
reservoir_weight[157][81],
reservoir_weight[157][82],
reservoir_weight[157][83],
reservoir_weight[157][84],
reservoir_weight[157][85],
reservoir_weight[157][86],
reservoir_weight[157][87],
reservoir_weight[157][88],
reservoir_weight[157][89],
reservoir_weight[157][90],
reservoir_weight[157][91],
reservoir_weight[157][92],
reservoir_weight[157][93],
reservoir_weight[157][94],
reservoir_weight[157][95],
reservoir_weight[157][96],
reservoir_weight[157][97],
reservoir_weight[157][98],
reservoir_weight[157][99],
reservoir_weight[157][100],
reservoir_weight[157][101],
reservoir_weight[157][102],
reservoir_weight[157][103],
reservoir_weight[157][104],
reservoir_weight[157][105],
reservoir_weight[157][106],
reservoir_weight[157][107],
reservoir_weight[157][108],
reservoir_weight[157][109],
reservoir_weight[157][110],
reservoir_weight[157][111],
reservoir_weight[157][112],
reservoir_weight[157][113],
reservoir_weight[157][114],
reservoir_weight[157][115],
reservoir_weight[157][116],
reservoir_weight[157][117],
reservoir_weight[157][118],
reservoir_weight[157][119],
reservoir_weight[157][120],
reservoir_weight[157][121],
reservoir_weight[157][122],
reservoir_weight[157][123],
reservoir_weight[157][124],
reservoir_weight[157][125],
reservoir_weight[157][126],
reservoir_weight[157][127],
reservoir_weight[157][128],
reservoir_weight[157][129],
reservoir_weight[157][130],
reservoir_weight[157][131],
reservoir_weight[157][132],
reservoir_weight[157][133],
reservoir_weight[157][134],
reservoir_weight[157][135],
reservoir_weight[157][136],
reservoir_weight[157][137],
reservoir_weight[157][138],
reservoir_weight[157][139],
reservoir_weight[157][140],
reservoir_weight[157][141],
reservoir_weight[157][142],
reservoir_weight[157][143],
reservoir_weight[157][144],
reservoir_weight[157][145],
reservoir_weight[157][146],
reservoir_weight[157][147],
reservoir_weight[157][148],
reservoir_weight[157][149],
reservoir_weight[157][150],
reservoir_weight[157][151],
reservoir_weight[157][152],
reservoir_weight[157][153],
reservoir_weight[157][154],
reservoir_weight[157][155],
reservoir_weight[157][156],
reservoir_weight[157][157],
reservoir_weight[157][158],
reservoir_weight[157][159],
reservoir_weight[157][160],
reservoir_weight[157][161],
reservoir_weight[157][162],
reservoir_weight[157][163],
reservoir_weight[157][164],
reservoir_weight[157][165],
reservoir_weight[157][166],
reservoir_weight[157][167],
reservoir_weight[157][168],
reservoir_weight[157][169],
reservoir_weight[157][170],
reservoir_weight[157][171],
reservoir_weight[157][172],
reservoir_weight[157][173],
reservoir_weight[157][174],
reservoir_weight[157][175],
reservoir_weight[157][176],
reservoir_weight[157][177],
reservoir_weight[157][178],
reservoir_weight[157][179],
reservoir_weight[157][180],
reservoir_weight[157][181],
reservoir_weight[157][182],
reservoir_weight[157][183],
reservoir_weight[157][184],
reservoir_weight[157][185],
reservoir_weight[157][186],
reservoir_weight[157][187],
reservoir_weight[157][188],
reservoir_weight[157][189],
reservoir_weight[157][190],
reservoir_weight[157][191],
reservoir_weight[157][192],
reservoir_weight[157][193],
reservoir_weight[157][194],
reservoir_weight[157][195],
reservoir_weight[157][196],
reservoir_weight[157][197],
reservoir_weight[157][198],
reservoir_weight[157][199]
},
{reservoir_weight[158][0],
reservoir_weight[158][1],
reservoir_weight[158][2],
reservoir_weight[158][3],
reservoir_weight[158][4],
reservoir_weight[158][5],
reservoir_weight[158][6],
reservoir_weight[158][7],
reservoir_weight[158][8],
reservoir_weight[158][9],
reservoir_weight[158][10],
reservoir_weight[158][11],
reservoir_weight[158][12],
reservoir_weight[158][13],
reservoir_weight[158][14],
reservoir_weight[158][15],
reservoir_weight[158][16],
reservoir_weight[158][17],
reservoir_weight[158][18],
reservoir_weight[158][19],
reservoir_weight[158][20],
reservoir_weight[158][21],
reservoir_weight[158][22],
reservoir_weight[158][23],
reservoir_weight[158][24],
reservoir_weight[158][25],
reservoir_weight[158][26],
reservoir_weight[158][27],
reservoir_weight[158][28],
reservoir_weight[158][29],
reservoir_weight[158][30],
reservoir_weight[158][31],
reservoir_weight[158][32],
reservoir_weight[158][33],
reservoir_weight[158][34],
reservoir_weight[158][35],
reservoir_weight[158][36],
reservoir_weight[158][37],
reservoir_weight[158][38],
reservoir_weight[158][39],
reservoir_weight[158][40],
reservoir_weight[158][41],
reservoir_weight[158][42],
reservoir_weight[158][43],
reservoir_weight[158][44],
reservoir_weight[158][45],
reservoir_weight[158][46],
reservoir_weight[158][47],
reservoir_weight[158][48],
reservoir_weight[158][49],
reservoir_weight[158][50],
reservoir_weight[158][51],
reservoir_weight[158][52],
reservoir_weight[158][53],
reservoir_weight[158][54],
reservoir_weight[158][55],
reservoir_weight[158][56],
reservoir_weight[158][57],
reservoir_weight[158][58],
reservoir_weight[158][59],
reservoir_weight[158][60],
reservoir_weight[158][61],
reservoir_weight[158][62],
reservoir_weight[158][63],
reservoir_weight[158][64],
reservoir_weight[158][65],
reservoir_weight[158][66],
reservoir_weight[158][67],
reservoir_weight[158][68],
reservoir_weight[158][69],
reservoir_weight[158][70],
reservoir_weight[158][71],
reservoir_weight[158][72],
reservoir_weight[158][73],
reservoir_weight[158][74],
reservoir_weight[158][75],
reservoir_weight[158][76],
reservoir_weight[158][77],
reservoir_weight[158][78],
reservoir_weight[158][79],
reservoir_weight[158][80],
reservoir_weight[158][81],
reservoir_weight[158][82],
reservoir_weight[158][83],
reservoir_weight[158][84],
reservoir_weight[158][85],
reservoir_weight[158][86],
reservoir_weight[158][87],
reservoir_weight[158][88],
reservoir_weight[158][89],
reservoir_weight[158][90],
reservoir_weight[158][91],
reservoir_weight[158][92],
reservoir_weight[158][93],
reservoir_weight[158][94],
reservoir_weight[158][95],
reservoir_weight[158][96],
reservoir_weight[158][97],
reservoir_weight[158][98],
reservoir_weight[158][99],
reservoir_weight[158][100],
reservoir_weight[158][101],
reservoir_weight[158][102],
reservoir_weight[158][103],
reservoir_weight[158][104],
reservoir_weight[158][105],
reservoir_weight[158][106],
reservoir_weight[158][107],
reservoir_weight[158][108],
reservoir_weight[158][109],
reservoir_weight[158][110],
reservoir_weight[158][111],
reservoir_weight[158][112],
reservoir_weight[158][113],
reservoir_weight[158][114],
reservoir_weight[158][115],
reservoir_weight[158][116],
reservoir_weight[158][117],
reservoir_weight[158][118],
reservoir_weight[158][119],
reservoir_weight[158][120],
reservoir_weight[158][121],
reservoir_weight[158][122],
reservoir_weight[158][123],
reservoir_weight[158][124],
reservoir_weight[158][125],
reservoir_weight[158][126],
reservoir_weight[158][127],
reservoir_weight[158][128],
reservoir_weight[158][129],
reservoir_weight[158][130],
reservoir_weight[158][131],
reservoir_weight[158][132],
reservoir_weight[158][133],
reservoir_weight[158][134],
reservoir_weight[158][135],
reservoir_weight[158][136],
reservoir_weight[158][137],
reservoir_weight[158][138],
reservoir_weight[158][139],
reservoir_weight[158][140],
reservoir_weight[158][141],
reservoir_weight[158][142],
reservoir_weight[158][143],
reservoir_weight[158][144],
reservoir_weight[158][145],
reservoir_weight[158][146],
reservoir_weight[158][147],
reservoir_weight[158][148],
reservoir_weight[158][149],
reservoir_weight[158][150],
reservoir_weight[158][151],
reservoir_weight[158][152],
reservoir_weight[158][153],
reservoir_weight[158][154],
reservoir_weight[158][155],
reservoir_weight[158][156],
reservoir_weight[158][157],
reservoir_weight[158][158],
reservoir_weight[158][159],
reservoir_weight[158][160],
reservoir_weight[158][161],
reservoir_weight[158][162],
reservoir_weight[158][163],
reservoir_weight[158][164],
reservoir_weight[158][165],
reservoir_weight[158][166],
reservoir_weight[158][167],
reservoir_weight[158][168],
reservoir_weight[158][169],
reservoir_weight[158][170],
reservoir_weight[158][171],
reservoir_weight[158][172],
reservoir_weight[158][173],
reservoir_weight[158][174],
reservoir_weight[158][175],
reservoir_weight[158][176],
reservoir_weight[158][177],
reservoir_weight[158][178],
reservoir_weight[158][179],
reservoir_weight[158][180],
reservoir_weight[158][181],
reservoir_weight[158][182],
reservoir_weight[158][183],
reservoir_weight[158][184],
reservoir_weight[158][185],
reservoir_weight[158][186],
reservoir_weight[158][187],
reservoir_weight[158][188],
reservoir_weight[158][189],
reservoir_weight[158][190],
reservoir_weight[158][191],
reservoir_weight[158][192],
reservoir_weight[158][193],
reservoir_weight[158][194],
reservoir_weight[158][195],
reservoir_weight[158][196],
reservoir_weight[158][197],
reservoir_weight[158][198],
reservoir_weight[158][199]
},
{reservoir_weight[159][0],
reservoir_weight[159][1],
reservoir_weight[159][2],
reservoir_weight[159][3],
reservoir_weight[159][4],
reservoir_weight[159][5],
reservoir_weight[159][6],
reservoir_weight[159][7],
reservoir_weight[159][8],
reservoir_weight[159][9],
reservoir_weight[159][10],
reservoir_weight[159][11],
reservoir_weight[159][12],
reservoir_weight[159][13],
reservoir_weight[159][14],
reservoir_weight[159][15],
reservoir_weight[159][16],
reservoir_weight[159][17],
reservoir_weight[159][18],
reservoir_weight[159][19],
reservoir_weight[159][20],
reservoir_weight[159][21],
reservoir_weight[159][22],
reservoir_weight[159][23],
reservoir_weight[159][24],
reservoir_weight[159][25],
reservoir_weight[159][26],
reservoir_weight[159][27],
reservoir_weight[159][28],
reservoir_weight[159][29],
reservoir_weight[159][30],
reservoir_weight[159][31],
reservoir_weight[159][32],
reservoir_weight[159][33],
reservoir_weight[159][34],
reservoir_weight[159][35],
reservoir_weight[159][36],
reservoir_weight[159][37],
reservoir_weight[159][38],
reservoir_weight[159][39],
reservoir_weight[159][40],
reservoir_weight[159][41],
reservoir_weight[159][42],
reservoir_weight[159][43],
reservoir_weight[159][44],
reservoir_weight[159][45],
reservoir_weight[159][46],
reservoir_weight[159][47],
reservoir_weight[159][48],
reservoir_weight[159][49],
reservoir_weight[159][50],
reservoir_weight[159][51],
reservoir_weight[159][52],
reservoir_weight[159][53],
reservoir_weight[159][54],
reservoir_weight[159][55],
reservoir_weight[159][56],
reservoir_weight[159][57],
reservoir_weight[159][58],
reservoir_weight[159][59],
reservoir_weight[159][60],
reservoir_weight[159][61],
reservoir_weight[159][62],
reservoir_weight[159][63],
reservoir_weight[159][64],
reservoir_weight[159][65],
reservoir_weight[159][66],
reservoir_weight[159][67],
reservoir_weight[159][68],
reservoir_weight[159][69],
reservoir_weight[159][70],
reservoir_weight[159][71],
reservoir_weight[159][72],
reservoir_weight[159][73],
reservoir_weight[159][74],
reservoir_weight[159][75],
reservoir_weight[159][76],
reservoir_weight[159][77],
reservoir_weight[159][78],
reservoir_weight[159][79],
reservoir_weight[159][80],
reservoir_weight[159][81],
reservoir_weight[159][82],
reservoir_weight[159][83],
reservoir_weight[159][84],
reservoir_weight[159][85],
reservoir_weight[159][86],
reservoir_weight[159][87],
reservoir_weight[159][88],
reservoir_weight[159][89],
reservoir_weight[159][90],
reservoir_weight[159][91],
reservoir_weight[159][92],
reservoir_weight[159][93],
reservoir_weight[159][94],
reservoir_weight[159][95],
reservoir_weight[159][96],
reservoir_weight[159][97],
reservoir_weight[159][98],
reservoir_weight[159][99],
reservoir_weight[159][100],
reservoir_weight[159][101],
reservoir_weight[159][102],
reservoir_weight[159][103],
reservoir_weight[159][104],
reservoir_weight[159][105],
reservoir_weight[159][106],
reservoir_weight[159][107],
reservoir_weight[159][108],
reservoir_weight[159][109],
reservoir_weight[159][110],
reservoir_weight[159][111],
reservoir_weight[159][112],
reservoir_weight[159][113],
reservoir_weight[159][114],
reservoir_weight[159][115],
reservoir_weight[159][116],
reservoir_weight[159][117],
reservoir_weight[159][118],
reservoir_weight[159][119],
reservoir_weight[159][120],
reservoir_weight[159][121],
reservoir_weight[159][122],
reservoir_weight[159][123],
reservoir_weight[159][124],
reservoir_weight[159][125],
reservoir_weight[159][126],
reservoir_weight[159][127],
reservoir_weight[159][128],
reservoir_weight[159][129],
reservoir_weight[159][130],
reservoir_weight[159][131],
reservoir_weight[159][132],
reservoir_weight[159][133],
reservoir_weight[159][134],
reservoir_weight[159][135],
reservoir_weight[159][136],
reservoir_weight[159][137],
reservoir_weight[159][138],
reservoir_weight[159][139],
reservoir_weight[159][140],
reservoir_weight[159][141],
reservoir_weight[159][142],
reservoir_weight[159][143],
reservoir_weight[159][144],
reservoir_weight[159][145],
reservoir_weight[159][146],
reservoir_weight[159][147],
reservoir_weight[159][148],
reservoir_weight[159][149],
reservoir_weight[159][150],
reservoir_weight[159][151],
reservoir_weight[159][152],
reservoir_weight[159][153],
reservoir_weight[159][154],
reservoir_weight[159][155],
reservoir_weight[159][156],
reservoir_weight[159][157],
reservoir_weight[159][158],
reservoir_weight[159][159],
reservoir_weight[159][160],
reservoir_weight[159][161],
reservoir_weight[159][162],
reservoir_weight[159][163],
reservoir_weight[159][164],
reservoir_weight[159][165],
reservoir_weight[159][166],
reservoir_weight[159][167],
reservoir_weight[159][168],
reservoir_weight[159][169],
reservoir_weight[159][170],
reservoir_weight[159][171],
reservoir_weight[159][172],
reservoir_weight[159][173],
reservoir_weight[159][174],
reservoir_weight[159][175],
reservoir_weight[159][176],
reservoir_weight[159][177],
reservoir_weight[159][178],
reservoir_weight[159][179],
reservoir_weight[159][180],
reservoir_weight[159][181],
reservoir_weight[159][182],
reservoir_weight[159][183],
reservoir_weight[159][184],
reservoir_weight[159][185],
reservoir_weight[159][186],
reservoir_weight[159][187],
reservoir_weight[159][188],
reservoir_weight[159][189],
reservoir_weight[159][190],
reservoir_weight[159][191],
reservoir_weight[159][192],
reservoir_weight[159][193],
reservoir_weight[159][194],
reservoir_weight[159][195],
reservoir_weight[159][196],
reservoir_weight[159][197],
reservoir_weight[159][198],
reservoir_weight[159][199]
},
{reservoir_weight[160][0],
reservoir_weight[160][1],
reservoir_weight[160][2],
reservoir_weight[160][3],
reservoir_weight[160][4],
reservoir_weight[160][5],
reservoir_weight[160][6],
reservoir_weight[160][7],
reservoir_weight[160][8],
reservoir_weight[160][9],
reservoir_weight[160][10],
reservoir_weight[160][11],
reservoir_weight[160][12],
reservoir_weight[160][13],
reservoir_weight[160][14],
reservoir_weight[160][15],
reservoir_weight[160][16],
reservoir_weight[160][17],
reservoir_weight[160][18],
reservoir_weight[160][19],
reservoir_weight[160][20],
reservoir_weight[160][21],
reservoir_weight[160][22],
reservoir_weight[160][23],
reservoir_weight[160][24],
reservoir_weight[160][25],
reservoir_weight[160][26],
reservoir_weight[160][27],
reservoir_weight[160][28],
reservoir_weight[160][29],
reservoir_weight[160][30],
reservoir_weight[160][31],
reservoir_weight[160][32],
reservoir_weight[160][33],
reservoir_weight[160][34],
reservoir_weight[160][35],
reservoir_weight[160][36],
reservoir_weight[160][37],
reservoir_weight[160][38],
reservoir_weight[160][39],
reservoir_weight[160][40],
reservoir_weight[160][41],
reservoir_weight[160][42],
reservoir_weight[160][43],
reservoir_weight[160][44],
reservoir_weight[160][45],
reservoir_weight[160][46],
reservoir_weight[160][47],
reservoir_weight[160][48],
reservoir_weight[160][49],
reservoir_weight[160][50],
reservoir_weight[160][51],
reservoir_weight[160][52],
reservoir_weight[160][53],
reservoir_weight[160][54],
reservoir_weight[160][55],
reservoir_weight[160][56],
reservoir_weight[160][57],
reservoir_weight[160][58],
reservoir_weight[160][59],
reservoir_weight[160][60],
reservoir_weight[160][61],
reservoir_weight[160][62],
reservoir_weight[160][63],
reservoir_weight[160][64],
reservoir_weight[160][65],
reservoir_weight[160][66],
reservoir_weight[160][67],
reservoir_weight[160][68],
reservoir_weight[160][69],
reservoir_weight[160][70],
reservoir_weight[160][71],
reservoir_weight[160][72],
reservoir_weight[160][73],
reservoir_weight[160][74],
reservoir_weight[160][75],
reservoir_weight[160][76],
reservoir_weight[160][77],
reservoir_weight[160][78],
reservoir_weight[160][79],
reservoir_weight[160][80],
reservoir_weight[160][81],
reservoir_weight[160][82],
reservoir_weight[160][83],
reservoir_weight[160][84],
reservoir_weight[160][85],
reservoir_weight[160][86],
reservoir_weight[160][87],
reservoir_weight[160][88],
reservoir_weight[160][89],
reservoir_weight[160][90],
reservoir_weight[160][91],
reservoir_weight[160][92],
reservoir_weight[160][93],
reservoir_weight[160][94],
reservoir_weight[160][95],
reservoir_weight[160][96],
reservoir_weight[160][97],
reservoir_weight[160][98],
reservoir_weight[160][99],
reservoir_weight[160][100],
reservoir_weight[160][101],
reservoir_weight[160][102],
reservoir_weight[160][103],
reservoir_weight[160][104],
reservoir_weight[160][105],
reservoir_weight[160][106],
reservoir_weight[160][107],
reservoir_weight[160][108],
reservoir_weight[160][109],
reservoir_weight[160][110],
reservoir_weight[160][111],
reservoir_weight[160][112],
reservoir_weight[160][113],
reservoir_weight[160][114],
reservoir_weight[160][115],
reservoir_weight[160][116],
reservoir_weight[160][117],
reservoir_weight[160][118],
reservoir_weight[160][119],
reservoir_weight[160][120],
reservoir_weight[160][121],
reservoir_weight[160][122],
reservoir_weight[160][123],
reservoir_weight[160][124],
reservoir_weight[160][125],
reservoir_weight[160][126],
reservoir_weight[160][127],
reservoir_weight[160][128],
reservoir_weight[160][129],
reservoir_weight[160][130],
reservoir_weight[160][131],
reservoir_weight[160][132],
reservoir_weight[160][133],
reservoir_weight[160][134],
reservoir_weight[160][135],
reservoir_weight[160][136],
reservoir_weight[160][137],
reservoir_weight[160][138],
reservoir_weight[160][139],
reservoir_weight[160][140],
reservoir_weight[160][141],
reservoir_weight[160][142],
reservoir_weight[160][143],
reservoir_weight[160][144],
reservoir_weight[160][145],
reservoir_weight[160][146],
reservoir_weight[160][147],
reservoir_weight[160][148],
reservoir_weight[160][149],
reservoir_weight[160][150],
reservoir_weight[160][151],
reservoir_weight[160][152],
reservoir_weight[160][153],
reservoir_weight[160][154],
reservoir_weight[160][155],
reservoir_weight[160][156],
reservoir_weight[160][157],
reservoir_weight[160][158],
reservoir_weight[160][159],
reservoir_weight[160][160],
reservoir_weight[160][161],
reservoir_weight[160][162],
reservoir_weight[160][163],
reservoir_weight[160][164],
reservoir_weight[160][165],
reservoir_weight[160][166],
reservoir_weight[160][167],
reservoir_weight[160][168],
reservoir_weight[160][169],
reservoir_weight[160][170],
reservoir_weight[160][171],
reservoir_weight[160][172],
reservoir_weight[160][173],
reservoir_weight[160][174],
reservoir_weight[160][175],
reservoir_weight[160][176],
reservoir_weight[160][177],
reservoir_weight[160][178],
reservoir_weight[160][179],
reservoir_weight[160][180],
reservoir_weight[160][181],
reservoir_weight[160][182],
reservoir_weight[160][183],
reservoir_weight[160][184],
reservoir_weight[160][185],
reservoir_weight[160][186],
reservoir_weight[160][187],
reservoir_weight[160][188],
reservoir_weight[160][189],
reservoir_weight[160][190],
reservoir_weight[160][191],
reservoir_weight[160][192],
reservoir_weight[160][193],
reservoir_weight[160][194],
reservoir_weight[160][195],
reservoir_weight[160][196],
reservoir_weight[160][197],
reservoir_weight[160][198],
reservoir_weight[160][199]
},
{reservoir_weight[161][0],
reservoir_weight[161][1],
reservoir_weight[161][2],
reservoir_weight[161][3],
reservoir_weight[161][4],
reservoir_weight[161][5],
reservoir_weight[161][6],
reservoir_weight[161][7],
reservoir_weight[161][8],
reservoir_weight[161][9],
reservoir_weight[161][10],
reservoir_weight[161][11],
reservoir_weight[161][12],
reservoir_weight[161][13],
reservoir_weight[161][14],
reservoir_weight[161][15],
reservoir_weight[161][16],
reservoir_weight[161][17],
reservoir_weight[161][18],
reservoir_weight[161][19],
reservoir_weight[161][20],
reservoir_weight[161][21],
reservoir_weight[161][22],
reservoir_weight[161][23],
reservoir_weight[161][24],
reservoir_weight[161][25],
reservoir_weight[161][26],
reservoir_weight[161][27],
reservoir_weight[161][28],
reservoir_weight[161][29],
reservoir_weight[161][30],
reservoir_weight[161][31],
reservoir_weight[161][32],
reservoir_weight[161][33],
reservoir_weight[161][34],
reservoir_weight[161][35],
reservoir_weight[161][36],
reservoir_weight[161][37],
reservoir_weight[161][38],
reservoir_weight[161][39],
reservoir_weight[161][40],
reservoir_weight[161][41],
reservoir_weight[161][42],
reservoir_weight[161][43],
reservoir_weight[161][44],
reservoir_weight[161][45],
reservoir_weight[161][46],
reservoir_weight[161][47],
reservoir_weight[161][48],
reservoir_weight[161][49],
reservoir_weight[161][50],
reservoir_weight[161][51],
reservoir_weight[161][52],
reservoir_weight[161][53],
reservoir_weight[161][54],
reservoir_weight[161][55],
reservoir_weight[161][56],
reservoir_weight[161][57],
reservoir_weight[161][58],
reservoir_weight[161][59],
reservoir_weight[161][60],
reservoir_weight[161][61],
reservoir_weight[161][62],
reservoir_weight[161][63],
reservoir_weight[161][64],
reservoir_weight[161][65],
reservoir_weight[161][66],
reservoir_weight[161][67],
reservoir_weight[161][68],
reservoir_weight[161][69],
reservoir_weight[161][70],
reservoir_weight[161][71],
reservoir_weight[161][72],
reservoir_weight[161][73],
reservoir_weight[161][74],
reservoir_weight[161][75],
reservoir_weight[161][76],
reservoir_weight[161][77],
reservoir_weight[161][78],
reservoir_weight[161][79],
reservoir_weight[161][80],
reservoir_weight[161][81],
reservoir_weight[161][82],
reservoir_weight[161][83],
reservoir_weight[161][84],
reservoir_weight[161][85],
reservoir_weight[161][86],
reservoir_weight[161][87],
reservoir_weight[161][88],
reservoir_weight[161][89],
reservoir_weight[161][90],
reservoir_weight[161][91],
reservoir_weight[161][92],
reservoir_weight[161][93],
reservoir_weight[161][94],
reservoir_weight[161][95],
reservoir_weight[161][96],
reservoir_weight[161][97],
reservoir_weight[161][98],
reservoir_weight[161][99],
reservoir_weight[161][100],
reservoir_weight[161][101],
reservoir_weight[161][102],
reservoir_weight[161][103],
reservoir_weight[161][104],
reservoir_weight[161][105],
reservoir_weight[161][106],
reservoir_weight[161][107],
reservoir_weight[161][108],
reservoir_weight[161][109],
reservoir_weight[161][110],
reservoir_weight[161][111],
reservoir_weight[161][112],
reservoir_weight[161][113],
reservoir_weight[161][114],
reservoir_weight[161][115],
reservoir_weight[161][116],
reservoir_weight[161][117],
reservoir_weight[161][118],
reservoir_weight[161][119],
reservoir_weight[161][120],
reservoir_weight[161][121],
reservoir_weight[161][122],
reservoir_weight[161][123],
reservoir_weight[161][124],
reservoir_weight[161][125],
reservoir_weight[161][126],
reservoir_weight[161][127],
reservoir_weight[161][128],
reservoir_weight[161][129],
reservoir_weight[161][130],
reservoir_weight[161][131],
reservoir_weight[161][132],
reservoir_weight[161][133],
reservoir_weight[161][134],
reservoir_weight[161][135],
reservoir_weight[161][136],
reservoir_weight[161][137],
reservoir_weight[161][138],
reservoir_weight[161][139],
reservoir_weight[161][140],
reservoir_weight[161][141],
reservoir_weight[161][142],
reservoir_weight[161][143],
reservoir_weight[161][144],
reservoir_weight[161][145],
reservoir_weight[161][146],
reservoir_weight[161][147],
reservoir_weight[161][148],
reservoir_weight[161][149],
reservoir_weight[161][150],
reservoir_weight[161][151],
reservoir_weight[161][152],
reservoir_weight[161][153],
reservoir_weight[161][154],
reservoir_weight[161][155],
reservoir_weight[161][156],
reservoir_weight[161][157],
reservoir_weight[161][158],
reservoir_weight[161][159],
reservoir_weight[161][160],
reservoir_weight[161][161],
reservoir_weight[161][162],
reservoir_weight[161][163],
reservoir_weight[161][164],
reservoir_weight[161][165],
reservoir_weight[161][166],
reservoir_weight[161][167],
reservoir_weight[161][168],
reservoir_weight[161][169],
reservoir_weight[161][170],
reservoir_weight[161][171],
reservoir_weight[161][172],
reservoir_weight[161][173],
reservoir_weight[161][174],
reservoir_weight[161][175],
reservoir_weight[161][176],
reservoir_weight[161][177],
reservoir_weight[161][178],
reservoir_weight[161][179],
reservoir_weight[161][180],
reservoir_weight[161][181],
reservoir_weight[161][182],
reservoir_weight[161][183],
reservoir_weight[161][184],
reservoir_weight[161][185],
reservoir_weight[161][186],
reservoir_weight[161][187],
reservoir_weight[161][188],
reservoir_weight[161][189],
reservoir_weight[161][190],
reservoir_weight[161][191],
reservoir_weight[161][192],
reservoir_weight[161][193],
reservoir_weight[161][194],
reservoir_weight[161][195],
reservoir_weight[161][196],
reservoir_weight[161][197],
reservoir_weight[161][198],
reservoir_weight[161][199]
},
{reservoir_weight[162][0],
reservoir_weight[162][1],
reservoir_weight[162][2],
reservoir_weight[162][3],
reservoir_weight[162][4],
reservoir_weight[162][5],
reservoir_weight[162][6],
reservoir_weight[162][7],
reservoir_weight[162][8],
reservoir_weight[162][9],
reservoir_weight[162][10],
reservoir_weight[162][11],
reservoir_weight[162][12],
reservoir_weight[162][13],
reservoir_weight[162][14],
reservoir_weight[162][15],
reservoir_weight[162][16],
reservoir_weight[162][17],
reservoir_weight[162][18],
reservoir_weight[162][19],
reservoir_weight[162][20],
reservoir_weight[162][21],
reservoir_weight[162][22],
reservoir_weight[162][23],
reservoir_weight[162][24],
reservoir_weight[162][25],
reservoir_weight[162][26],
reservoir_weight[162][27],
reservoir_weight[162][28],
reservoir_weight[162][29],
reservoir_weight[162][30],
reservoir_weight[162][31],
reservoir_weight[162][32],
reservoir_weight[162][33],
reservoir_weight[162][34],
reservoir_weight[162][35],
reservoir_weight[162][36],
reservoir_weight[162][37],
reservoir_weight[162][38],
reservoir_weight[162][39],
reservoir_weight[162][40],
reservoir_weight[162][41],
reservoir_weight[162][42],
reservoir_weight[162][43],
reservoir_weight[162][44],
reservoir_weight[162][45],
reservoir_weight[162][46],
reservoir_weight[162][47],
reservoir_weight[162][48],
reservoir_weight[162][49],
reservoir_weight[162][50],
reservoir_weight[162][51],
reservoir_weight[162][52],
reservoir_weight[162][53],
reservoir_weight[162][54],
reservoir_weight[162][55],
reservoir_weight[162][56],
reservoir_weight[162][57],
reservoir_weight[162][58],
reservoir_weight[162][59],
reservoir_weight[162][60],
reservoir_weight[162][61],
reservoir_weight[162][62],
reservoir_weight[162][63],
reservoir_weight[162][64],
reservoir_weight[162][65],
reservoir_weight[162][66],
reservoir_weight[162][67],
reservoir_weight[162][68],
reservoir_weight[162][69],
reservoir_weight[162][70],
reservoir_weight[162][71],
reservoir_weight[162][72],
reservoir_weight[162][73],
reservoir_weight[162][74],
reservoir_weight[162][75],
reservoir_weight[162][76],
reservoir_weight[162][77],
reservoir_weight[162][78],
reservoir_weight[162][79],
reservoir_weight[162][80],
reservoir_weight[162][81],
reservoir_weight[162][82],
reservoir_weight[162][83],
reservoir_weight[162][84],
reservoir_weight[162][85],
reservoir_weight[162][86],
reservoir_weight[162][87],
reservoir_weight[162][88],
reservoir_weight[162][89],
reservoir_weight[162][90],
reservoir_weight[162][91],
reservoir_weight[162][92],
reservoir_weight[162][93],
reservoir_weight[162][94],
reservoir_weight[162][95],
reservoir_weight[162][96],
reservoir_weight[162][97],
reservoir_weight[162][98],
reservoir_weight[162][99],
reservoir_weight[162][100],
reservoir_weight[162][101],
reservoir_weight[162][102],
reservoir_weight[162][103],
reservoir_weight[162][104],
reservoir_weight[162][105],
reservoir_weight[162][106],
reservoir_weight[162][107],
reservoir_weight[162][108],
reservoir_weight[162][109],
reservoir_weight[162][110],
reservoir_weight[162][111],
reservoir_weight[162][112],
reservoir_weight[162][113],
reservoir_weight[162][114],
reservoir_weight[162][115],
reservoir_weight[162][116],
reservoir_weight[162][117],
reservoir_weight[162][118],
reservoir_weight[162][119],
reservoir_weight[162][120],
reservoir_weight[162][121],
reservoir_weight[162][122],
reservoir_weight[162][123],
reservoir_weight[162][124],
reservoir_weight[162][125],
reservoir_weight[162][126],
reservoir_weight[162][127],
reservoir_weight[162][128],
reservoir_weight[162][129],
reservoir_weight[162][130],
reservoir_weight[162][131],
reservoir_weight[162][132],
reservoir_weight[162][133],
reservoir_weight[162][134],
reservoir_weight[162][135],
reservoir_weight[162][136],
reservoir_weight[162][137],
reservoir_weight[162][138],
reservoir_weight[162][139],
reservoir_weight[162][140],
reservoir_weight[162][141],
reservoir_weight[162][142],
reservoir_weight[162][143],
reservoir_weight[162][144],
reservoir_weight[162][145],
reservoir_weight[162][146],
reservoir_weight[162][147],
reservoir_weight[162][148],
reservoir_weight[162][149],
reservoir_weight[162][150],
reservoir_weight[162][151],
reservoir_weight[162][152],
reservoir_weight[162][153],
reservoir_weight[162][154],
reservoir_weight[162][155],
reservoir_weight[162][156],
reservoir_weight[162][157],
reservoir_weight[162][158],
reservoir_weight[162][159],
reservoir_weight[162][160],
reservoir_weight[162][161],
reservoir_weight[162][162],
reservoir_weight[162][163],
reservoir_weight[162][164],
reservoir_weight[162][165],
reservoir_weight[162][166],
reservoir_weight[162][167],
reservoir_weight[162][168],
reservoir_weight[162][169],
reservoir_weight[162][170],
reservoir_weight[162][171],
reservoir_weight[162][172],
reservoir_weight[162][173],
reservoir_weight[162][174],
reservoir_weight[162][175],
reservoir_weight[162][176],
reservoir_weight[162][177],
reservoir_weight[162][178],
reservoir_weight[162][179],
reservoir_weight[162][180],
reservoir_weight[162][181],
reservoir_weight[162][182],
reservoir_weight[162][183],
reservoir_weight[162][184],
reservoir_weight[162][185],
reservoir_weight[162][186],
reservoir_weight[162][187],
reservoir_weight[162][188],
reservoir_weight[162][189],
reservoir_weight[162][190],
reservoir_weight[162][191],
reservoir_weight[162][192],
reservoir_weight[162][193],
reservoir_weight[162][194],
reservoir_weight[162][195],
reservoir_weight[162][196],
reservoir_weight[162][197],
reservoir_weight[162][198],
reservoir_weight[162][199]
},
{reservoir_weight[163][0],
reservoir_weight[163][1],
reservoir_weight[163][2],
reservoir_weight[163][3],
reservoir_weight[163][4],
reservoir_weight[163][5],
reservoir_weight[163][6],
reservoir_weight[163][7],
reservoir_weight[163][8],
reservoir_weight[163][9],
reservoir_weight[163][10],
reservoir_weight[163][11],
reservoir_weight[163][12],
reservoir_weight[163][13],
reservoir_weight[163][14],
reservoir_weight[163][15],
reservoir_weight[163][16],
reservoir_weight[163][17],
reservoir_weight[163][18],
reservoir_weight[163][19],
reservoir_weight[163][20],
reservoir_weight[163][21],
reservoir_weight[163][22],
reservoir_weight[163][23],
reservoir_weight[163][24],
reservoir_weight[163][25],
reservoir_weight[163][26],
reservoir_weight[163][27],
reservoir_weight[163][28],
reservoir_weight[163][29],
reservoir_weight[163][30],
reservoir_weight[163][31],
reservoir_weight[163][32],
reservoir_weight[163][33],
reservoir_weight[163][34],
reservoir_weight[163][35],
reservoir_weight[163][36],
reservoir_weight[163][37],
reservoir_weight[163][38],
reservoir_weight[163][39],
reservoir_weight[163][40],
reservoir_weight[163][41],
reservoir_weight[163][42],
reservoir_weight[163][43],
reservoir_weight[163][44],
reservoir_weight[163][45],
reservoir_weight[163][46],
reservoir_weight[163][47],
reservoir_weight[163][48],
reservoir_weight[163][49],
reservoir_weight[163][50],
reservoir_weight[163][51],
reservoir_weight[163][52],
reservoir_weight[163][53],
reservoir_weight[163][54],
reservoir_weight[163][55],
reservoir_weight[163][56],
reservoir_weight[163][57],
reservoir_weight[163][58],
reservoir_weight[163][59],
reservoir_weight[163][60],
reservoir_weight[163][61],
reservoir_weight[163][62],
reservoir_weight[163][63],
reservoir_weight[163][64],
reservoir_weight[163][65],
reservoir_weight[163][66],
reservoir_weight[163][67],
reservoir_weight[163][68],
reservoir_weight[163][69],
reservoir_weight[163][70],
reservoir_weight[163][71],
reservoir_weight[163][72],
reservoir_weight[163][73],
reservoir_weight[163][74],
reservoir_weight[163][75],
reservoir_weight[163][76],
reservoir_weight[163][77],
reservoir_weight[163][78],
reservoir_weight[163][79],
reservoir_weight[163][80],
reservoir_weight[163][81],
reservoir_weight[163][82],
reservoir_weight[163][83],
reservoir_weight[163][84],
reservoir_weight[163][85],
reservoir_weight[163][86],
reservoir_weight[163][87],
reservoir_weight[163][88],
reservoir_weight[163][89],
reservoir_weight[163][90],
reservoir_weight[163][91],
reservoir_weight[163][92],
reservoir_weight[163][93],
reservoir_weight[163][94],
reservoir_weight[163][95],
reservoir_weight[163][96],
reservoir_weight[163][97],
reservoir_weight[163][98],
reservoir_weight[163][99],
reservoir_weight[163][100],
reservoir_weight[163][101],
reservoir_weight[163][102],
reservoir_weight[163][103],
reservoir_weight[163][104],
reservoir_weight[163][105],
reservoir_weight[163][106],
reservoir_weight[163][107],
reservoir_weight[163][108],
reservoir_weight[163][109],
reservoir_weight[163][110],
reservoir_weight[163][111],
reservoir_weight[163][112],
reservoir_weight[163][113],
reservoir_weight[163][114],
reservoir_weight[163][115],
reservoir_weight[163][116],
reservoir_weight[163][117],
reservoir_weight[163][118],
reservoir_weight[163][119],
reservoir_weight[163][120],
reservoir_weight[163][121],
reservoir_weight[163][122],
reservoir_weight[163][123],
reservoir_weight[163][124],
reservoir_weight[163][125],
reservoir_weight[163][126],
reservoir_weight[163][127],
reservoir_weight[163][128],
reservoir_weight[163][129],
reservoir_weight[163][130],
reservoir_weight[163][131],
reservoir_weight[163][132],
reservoir_weight[163][133],
reservoir_weight[163][134],
reservoir_weight[163][135],
reservoir_weight[163][136],
reservoir_weight[163][137],
reservoir_weight[163][138],
reservoir_weight[163][139],
reservoir_weight[163][140],
reservoir_weight[163][141],
reservoir_weight[163][142],
reservoir_weight[163][143],
reservoir_weight[163][144],
reservoir_weight[163][145],
reservoir_weight[163][146],
reservoir_weight[163][147],
reservoir_weight[163][148],
reservoir_weight[163][149],
reservoir_weight[163][150],
reservoir_weight[163][151],
reservoir_weight[163][152],
reservoir_weight[163][153],
reservoir_weight[163][154],
reservoir_weight[163][155],
reservoir_weight[163][156],
reservoir_weight[163][157],
reservoir_weight[163][158],
reservoir_weight[163][159],
reservoir_weight[163][160],
reservoir_weight[163][161],
reservoir_weight[163][162],
reservoir_weight[163][163],
reservoir_weight[163][164],
reservoir_weight[163][165],
reservoir_weight[163][166],
reservoir_weight[163][167],
reservoir_weight[163][168],
reservoir_weight[163][169],
reservoir_weight[163][170],
reservoir_weight[163][171],
reservoir_weight[163][172],
reservoir_weight[163][173],
reservoir_weight[163][174],
reservoir_weight[163][175],
reservoir_weight[163][176],
reservoir_weight[163][177],
reservoir_weight[163][178],
reservoir_weight[163][179],
reservoir_weight[163][180],
reservoir_weight[163][181],
reservoir_weight[163][182],
reservoir_weight[163][183],
reservoir_weight[163][184],
reservoir_weight[163][185],
reservoir_weight[163][186],
reservoir_weight[163][187],
reservoir_weight[163][188],
reservoir_weight[163][189],
reservoir_weight[163][190],
reservoir_weight[163][191],
reservoir_weight[163][192],
reservoir_weight[163][193],
reservoir_weight[163][194],
reservoir_weight[163][195],
reservoir_weight[163][196],
reservoir_weight[163][197],
reservoir_weight[163][198],
reservoir_weight[163][199]
},
{reservoir_weight[164][0],
reservoir_weight[164][1],
reservoir_weight[164][2],
reservoir_weight[164][3],
reservoir_weight[164][4],
reservoir_weight[164][5],
reservoir_weight[164][6],
reservoir_weight[164][7],
reservoir_weight[164][8],
reservoir_weight[164][9],
reservoir_weight[164][10],
reservoir_weight[164][11],
reservoir_weight[164][12],
reservoir_weight[164][13],
reservoir_weight[164][14],
reservoir_weight[164][15],
reservoir_weight[164][16],
reservoir_weight[164][17],
reservoir_weight[164][18],
reservoir_weight[164][19],
reservoir_weight[164][20],
reservoir_weight[164][21],
reservoir_weight[164][22],
reservoir_weight[164][23],
reservoir_weight[164][24],
reservoir_weight[164][25],
reservoir_weight[164][26],
reservoir_weight[164][27],
reservoir_weight[164][28],
reservoir_weight[164][29],
reservoir_weight[164][30],
reservoir_weight[164][31],
reservoir_weight[164][32],
reservoir_weight[164][33],
reservoir_weight[164][34],
reservoir_weight[164][35],
reservoir_weight[164][36],
reservoir_weight[164][37],
reservoir_weight[164][38],
reservoir_weight[164][39],
reservoir_weight[164][40],
reservoir_weight[164][41],
reservoir_weight[164][42],
reservoir_weight[164][43],
reservoir_weight[164][44],
reservoir_weight[164][45],
reservoir_weight[164][46],
reservoir_weight[164][47],
reservoir_weight[164][48],
reservoir_weight[164][49],
reservoir_weight[164][50],
reservoir_weight[164][51],
reservoir_weight[164][52],
reservoir_weight[164][53],
reservoir_weight[164][54],
reservoir_weight[164][55],
reservoir_weight[164][56],
reservoir_weight[164][57],
reservoir_weight[164][58],
reservoir_weight[164][59],
reservoir_weight[164][60],
reservoir_weight[164][61],
reservoir_weight[164][62],
reservoir_weight[164][63],
reservoir_weight[164][64],
reservoir_weight[164][65],
reservoir_weight[164][66],
reservoir_weight[164][67],
reservoir_weight[164][68],
reservoir_weight[164][69],
reservoir_weight[164][70],
reservoir_weight[164][71],
reservoir_weight[164][72],
reservoir_weight[164][73],
reservoir_weight[164][74],
reservoir_weight[164][75],
reservoir_weight[164][76],
reservoir_weight[164][77],
reservoir_weight[164][78],
reservoir_weight[164][79],
reservoir_weight[164][80],
reservoir_weight[164][81],
reservoir_weight[164][82],
reservoir_weight[164][83],
reservoir_weight[164][84],
reservoir_weight[164][85],
reservoir_weight[164][86],
reservoir_weight[164][87],
reservoir_weight[164][88],
reservoir_weight[164][89],
reservoir_weight[164][90],
reservoir_weight[164][91],
reservoir_weight[164][92],
reservoir_weight[164][93],
reservoir_weight[164][94],
reservoir_weight[164][95],
reservoir_weight[164][96],
reservoir_weight[164][97],
reservoir_weight[164][98],
reservoir_weight[164][99],
reservoir_weight[164][100],
reservoir_weight[164][101],
reservoir_weight[164][102],
reservoir_weight[164][103],
reservoir_weight[164][104],
reservoir_weight[164][105],
reservoir_weight[164][106],
reservoir_weight[164][107],
reservoir_weight[164][108],
reservoir_weight[164][109],
reservoir_weight[164][110],
reservoir_weight[164][111],
reservoir_weight[164][112],
reservoir_weight[164][113],
reservoir_weight[164][114],
reservoir_weight[164][115],
reservoir_weight[164][116],
reservoir_weight[164][117],
reservoir_weight[164][118],
reservoir_weight[164][119],
reservoir_weight[164][120],
reservoir_weight[164][121],
reservoir_weight[164][122],
reservoir_weight[164][123],
reservoir_weight[164][124],
reservoir_weight[164][125],
reservoir_weight[164][126],
reservoir_weight[164][127],
reservoir_weight[164][128],
reservoir_weight[164][129],
reservoir_weight[164][130],
reservoir_weight[164][131],
reservoir_weight[164][132],
reservoir_weight[164][133],
reservoir_weight[164][134],
reservoir_weight[164][135],
reservoir_weight[164][136],
reservoir_weight[164][137],
reservoir_weight[164][138],
reservoir_weight[164][139],
reservoir_weight[164][140],
reservoir_weight[164][141],
reservoir_weight[164][142],
reservoir_weight[164][143],
reservoir_weight[164][144],
reservoir_weight[164][145],
reservoir_weight[164][146],
reservoir_weight[164][147],
reservoir_weight[164][148],
reservoir_weight[164][149],
reservoir_weight[164][150],
reservoir_weight[164][151],
reservoir_weight[164][152],
reservoir_weight[164][153],
reservoir_weight[164][154],
reservoir_weight[164][155],
reservoir_weight[164][156],
reservoir_weight[164][157],
reservoir_weight[164][158],
reservoir_weight[164][159],
reservoir_weight[164][160],
reservoir_weight[164][161],
reservoir_weight[164][162],
reservoir_weight[164][163],
reservoir_weight[164][164],
reservoir_weight[164][165],
reservoir_weight[164][166],
reservoir_weight[164][167],
reservoir_weight[164][168],
reservoir_weight[164][169],
reservoir_weight[164][170],
reservoir_weight[164][171],
reservoir_weight[164][172],
reservoir_weight[164][173],
reservoir_weight[164][174],
reservoir_weight[164][175],
reservoir_weight[164][176],
reservoir_weight[164][177],
reservoir_weight[164][178],
reservoir_weight[164][179],
reservoir_weight[164][180],
reservoir_weight[164][181],
reservoir_weight[164][182],
reservoir_weight[164][183],
reservoir_weight[164][184],
reservoir_weight[164][185],
reservoir_weight[164][186],
reservoir_weight[164][187],
reservoir_weight[164][188],
reservoir_weight[164][189],
reservoir_weight[164][190],
reservoir_weight[164][191],
reservoir_weight[164][192],
reservoir_weight[164][193],
reservoir_weight[164][194],
reservoir_weight[164][195],
reservoir_weight[164][196],
reservoir_weight[164][197],
reservoir_weight[164][198],
reservoir_weight[164][199]
},
{reservoir_weight[165][0],
reservoir_weight[165][1],
reservoir_weight[165][2],
reservoir_weight[165][3],
reservoir_weight[165][4],
reservoir_weight[165][5],
reservoir_weight[165][6],
reservoir_weight[165][7],
reservoir_weight[165][8],
reservoir_weight[165][9],
reservoir_weight[165][10],
reservoir_weight[165][11],
reservoir_weight[165][12],
reservoir_weight[165][13],
reservoir_weight[165][14],
reservoir_weight[165][15],
reservoir_weight[165][16],
reservoir_weight[165][17],
reservoir_weight[165][18],
reservoir_weight[165][19],
reservoir_weight[165][20],
reservoir_weight[165][21],
reservoir_weight[165][22],
reservoir_weight[165][23],
reservoir_weight[165][24],
reservoir_weight[165][25],
reservoir_weight[165][26],
reservoir_weight[165][27],
reservoir_weight[165][28],
reservoir_weight[165][29],
reservoir_weight[165][30],
reservoir_weight[165][31],
reservoir_weight[165][32],
reservoir_weight[165][33],
reservoir_weight[165][34],
reservoir_weight[165][35],
reservoir_weight[165][36],
reservoir_weight[165][37],
reservoir_weight[165][38],
reservoir_weight[165][39],
reservoir_weight[165][40],
reservoir_weight[165][41],
reservoir_weight[165][42],
reservoir_weight[165][43],
reservoir_weight[165][44],
reservoir_weight[165][45],
reservoir_weight[165][46],
reservoir_weight[165][47],
reservoir_weight[165][48],
reservoir_weight[165][49],
reservoir_weight[165][50],
reservoir_weight[165][51],
reservoir_weight[165][52],
reservoir_weight[165][53],
reservoir_weight[165][54],
reservoir_weight[165][55],
reservoir_weight[165][56],
reservoir_weight[165][57],
reservoir_weight[165][58],
reservoir_weight[165][59],
reservoir_weight[165][60],
reservoir_weight[165][61],
reservoir_weight[165][62],
reservoir_weight[165][63],
reservoir_weight[165][64],
reservoir_weight[165][65],
reservoir_weight[165][66],
reservoir_weight[165][67],
reservoir_weight[165][68],
reservoir_weight[165][69],
reservoir_weight[165][70],
reservoir_weight[165][71],
reservoir_weight[165][72],
reservoir_weight[165][73],
reservoir_weight[165][74],
reservoir_weight[165][75],
reservoir_weight[165][76],
reservoir_weight[165][77],
reservoir_weight[165][78],
reservoir_weight[165][79],
reservoir_weight[165][80],
reservoir_weight[165][81],
reservoir_weight[165][82],
reservoir_weight[165][83],
reservoir_weight[165][84],
reservoir_weight[165][85],
reservoir_weight[165][86],
reservoir_weight[165][87],
reservoir_weight[165][88],
reservoir_weight[165][89],
reservoir_weight[165][90],
reservoir_weight[165][91],
reservoir_weight[165][92],
reservoir_weight[165][93],
reservoir_weight[165][94],
reservoir_weight[165][95],
reservoir_weight[165][96],
reservoir_weight[165][97],
reservoir_weight[165][98],
reservoir_weight[165][99],
reservoir_weight[165][100],
reservoir_weight[165][101],
reservoir_weight[165][102],
reservoir_weight[165][103],
reservoir_weight[165][104],
reservoir_weight[165][105],
reservoir_weight[165][106],
reservoir_weight[165][107],
reservoir_weight[165][108],
reservoir_weight[165][109],
reservoir_weight[165][110],
reservoir_weight[165][111],
reservoir_weight[165][112],
reservoir_weight[165][113],
reservoir_weight[165][114],
reservoir_weight[165][115],
reservoir_weight[165][116],
reservoir_weight[165][117],
reservoir_weight[165][118],
reservoir_weight[165][119],
reservoir_weight[165][120],
reservoir_weight[165][121],
reservoir_weight[165][122],
reservoir_weight[165][123],
reservoir_weight[165][124],
reservoir_weight[165][125],
reservoir_weight[165][126],
reservoir_weight[165][127],
reservoir_weight[165][128],
reservoir_weight[165][129],
reservoir_weight[165][130],
reservoir_weight[165][131],
reservoir_weight[165][132],
reservoir_weight[165][133],
reservoir_weight[165][134],
reservoir_weight[165][135],
reservoir_weight[165][136],
reservoir_weight[165][137],
reservoir_weight[165][138],
reservoir_weight[165][139],
reservoir_weight[165][140],
reservoir_weight[165][141],
reservoir_weight[165][142],
reservoir_weight[165][143],
reservoir_weight[165][144],
reservoir_weight[165][145],
reservoir_weight[165][146],
reservoir_weight[165][147],
reservoir_weight[165][148],
reservoir_weight[165][149],
reservoir_weight[165][150],
reservoir_weight[165][151],
reservoir_weight[165][152],
reservoir_weight[165][153],
reservoir_weight[165][154],
reservoir_weight[165][155],
reservoir_weight[165][156],
reservoir_weight[165][157],
reservoir_weight[165][158],
reservoir_weight[165][159],
reservoir_weight[165][160],
reservoir_weight[165][161],
reservoir_weight[165][162],
reservoir_weight[165][163],
reservoir_weight[165][164],
reservoir_weight[165][165],
reservoir_weight[165][166],
reservoir_weight[165][167],
reservoir_weight[165][168],
reservoir_weight[165][169],
reservoir_weight[165][170],
reservoir_weight[165][171],
reservoir_weight[165][172],
reservoir_weight[165][173],
reservoir_weight[165][174],
reservoir_weight[165][175],
reservoir_weight[165][176],
reservoir_weight[165][177],
reservoir_weight[165][178],
reservoir_weight[165][179],
reservoir_weight[165][180],
reservoir_weight[165][181],
reservoir_weight[165][182],
reservoir_weight[165][183],
reservoir_weight[165][184],
reservoir_weight[165][185],
reservoir_weight[165][186],
reservoir_weight[165][187],
reservoir_weight[165][188],
reservoir_weight[165][189],
reservoir_weight[165][190],
reservoir_weight[165][191],
reservoir_weight[165][192],
reservoir_weight[165][193],
reservoir_weight[165][194],
reservoir_weight[165][195],
reservoir_weight[165][196],
reservoir_weight[165][197],
reservoir_weight[165][198],
reservoir_weight[165][199]
},
{reservoir_weight[166][0],
reservoir_weight[166][1],
reservoir_weight[166][2],
reservoir_weight[166][3],
reservoir_weight[166][4],
reservoir_weight[166][5],
reservoir_weight[166][6],
reservoir_weight[166][7],
reservoir_weight[166][8],
reservoir_weight[166][9],
reservoir_weight[166][10],
reservoir_weight[166][11],
reservoir_weight[166][12],
reservoir_weight[166][13],
reservoir_weight[166][14],
reservoir_weight[166][15],
reservoir_weight[166][16],
reservoir_weight[166][17],
reservoir_weight[166][18],
reservoir_weight[166][19],
reservoir_weight[166][20],
reservoir_weight[166][21],
reservoir_weight[166][22],
reservoir_weight[166][23],
reservoir_weight[166][24],
reservoir_weight[166][25],
reservoir_weight[166][26],
reservoir_weight[166][27],
reservoir_weight[166][28],
reservoir_weight[166][29],
reservoir_weight[166][30],
reservoir_weight[166][31],
reservoir_weight[166][32],
reservoir_weight[166][33],
reservoir_weight[166][34],
reservoir_weight[166][35],
reservoir_weight[166][36],
reservoir_weight[166][37],
reservoir_weight[166][38],
reservoir_weight[166][39],
reservoir_weight[166][40],
reservoir_weight[166][41],
reservoir_weight[166][42],
reservoir_weight[166][43],
reservoir_weight[166][44],
reservoir_weight[166][45],
reservoir_weight[166][46],
reservoir_weight[166][47],
reservoir_weight[166][48],
reservoir_weight[166][49],
reservoir_weight[166][50],
reservoir_weight[166][51],
reservoir_weight[166][52],
reservoir_weight[166][53],
reservoir_weight[166][54],
reservoir_weight[166][55],
reservoir_weight[166][56],
reservoir_weight[166][57],
reservoir_weight[166][58],
reservoir_weight[166][59],
reservoir_weight[166][60],
reservoir_weight[166][61],
reservoir_weight[166][62],
reservoir_weight[166][63],
reservoir_weight[166][64],
reservoir_weight[166][65],
reservoir_weight[166][66],
reservoir_weight[166][67],
reservoir_weight[166][68],
reservoir_weight[166][69],
reservoir_weight[166][70],
reservoir_weight[166][71],
reservoir_weight[166][72],
reservoir_weight[166][73],
reservoir_weight[166][74],
reservoir_weight[166][75],
reservoir_weight[166][76],
reservoir_weight[166][77],
reservoir_weight[166][78],
reservoir_weight[166][79],
reservoir_weight[166][80],
reservoir_weight[166][81],
reservoir_weight[166][82],
reservoir_weight[166][83],
reservoir_weight[166][84],
reservoir_weight[166][85],
reservoir_weight[166][86],
reservoir_weight[166][87],
reservoir_weight[166][88],
reservoir_weight[166][89],
reservoir_weight[166][90],
reservoir_weight[166][91],
reservoir_weight[166][92],
reservoir_weight[166][93],
reservoir_weight[166][94],
reservoir_weight[166][95],
reservoir_weight[166][96],
reservoir_weight[166][97],
reservoir_weight[166][98],
reservoir_weight[166][99],
reservoir_weight[166][100],
reservoir_weight[166][101],
reservoir_weight[166][102],
reservoir_weight[166][103],
reservoir_weight[166][104],
reservoir_weight[166][105],
reservoir_weight[166][106],
reservoir_weight[166][107],
reservoir_weight[166][108],
reservoir_weight[166][109],
reservoir_weight[166][110],
reservoir_weight[166][111],
reservoir_weight[166][112],
reservoir_weight[166][113],
reservoir_weight[166][114],
reservoir_weight[166][115],
reservoir_weight[166][116],
reservoir_weight[166][117],
reservoir_weight[166][118],
reservoir_weight[166][119],
reservoir_weight[166][120],
reservoir_weight[166][121],
reservoir_weight[166][122],
reservoir_weight[166][123],
reservoir_weight[166][124],
reservoir_weight[166][125],
reservoir_weight[166][126],
reservoir_weight[166][127],
reservoir_weight[166][128],
reservoir_weight[166][129],
reservoir_weight[166][130],
reservoir_weight[166][131],
reservoir_weight[166][132],
reservoir_weight[166][133],
reservoir_weight[166][134],
reservoir_weight[166][135],
reservoir_weight[166][136],
reservoir_weight[166][137],
reservoir_weight[166][138],
reservoir_weight[166][139],
reservoir_weight[166][140],
reservoir_weight[166][141],
reservoir_weight[166][142],
reservoir_weight[166][143],
reservoir_weight[166][144],
reservoir_weight[166][145],
reservoir_weight[166][146],
reservoir_weight[166][147],
reservoir_weight[166][148],
reservoir_weight[166][149],
reservoir_weight[166][150],
reservoir_weight[166][151],
reservoir_weight[166][152],
reservoir_weight[166][153],
reservoir_weight[166][154],
reservoir_weight[166][155],
reservoir_weight[166][156],
reservoir_weight[166][157],
reservoir_weight[166][158],
reservoir_weight[166][159],
reservoir_weight[166][160],
reservoir_weight[166][161],
reservoir_weight[166][162],
reservoir_weight[166][163],
reservoir_weight[166][164],
reservoir_weight[166][165],
reservoir_weight[166][166],
reservoir_weight[166][167],
reservoir_weight[166][168],
reservoir_weight[166][169],
reservoir_weight[166][170],
reservoir_weight[166][171],
reservoir_weight[166][172],
reservoir_weight[166][173],
reservoir_weight[166][174],
reservoir_weight[166][175],
reservoir_weight[166][176],
reservoir_weight[166][177],
reservoir_weight[166][178],
reservoir_weight[166][179],
reservoir_weight[166][180],
reservoir_weight[166][181],
reservoir_weight[166][182],
reservoir_weight[166][183],
reservoir_weight[166][184],
reservoir_weight[166][185],
reservoir_weight[166][186],
reservoir_weight[166][187],
reservoir_weight[166][188],
reservoir_weight[166][189],
reservoir_weight[166][190],
reservoir_weight[166][191],
reservoir_weight[166][192],
reservoir_weight[166][193],
reservoir_weight[166][194],
reservoir_weight[166][195],
reservoir_weight[166][196],
reservoir_weight[166][197],
reservoir_weight[166][198],
reservoir_weight[166][199]
},
{reservoir_weight[167][0],
reservoir_weight[167][1],
reservoir_weight[167][2],
reservoir_weight[167][3],
reservoir_weight[167][4],
reservoir_weight[167][5],
reservoir_weight[167][6],
reservoir_weight[167][7],
reservoir_weight[167][8],
reservoir_weight[167][9],
reservoir_weight[167][10],
reservoir_weight[167][11],
reservoir_weight[167][12],
reservoir_weight[167][13],
reservoir_weight[167][14],
reservoir_weight[167][15],
reservoir_weight[167][16],
reservoir_weight[167][17],
reservoir_weight[167][18],
reservoir_weight[167][19],
reservoir_weight[167][20],
reservoir_weight[167][21],
reservoir_weight[167][22],
reservoir_weight[167][23],
reservoir_weight[167][24],
reservoir_weight[167][25],
reservoir_weight[167][26],
reservoir_weight[167][27],
reservoir_weight[167][28],
reservoir_weight[167][29],
reservoir_weight[167][30],
reservoir_weight[167][31],
reservoir_weight[167][32],
reservoir_weight[167][33],
reservoir_weight[167][34],
reservoir_weight[167][35],
reservoir_weight[167][36],
reservoir_weight[167][37],
reservoir_weight[167][38],
reservoir_weight[167][39],
reservoir_weight[167][40],
reservoir_weight[167][41],
reservoir_weight[167][42],
reservoir_weight[167][43],
reservoir_weight[167][44],
reservoir_weight[167][45],
reservoir_weight[167][46],
reservoir_weight[167][47],
reservoir_weight[167][48],
reservoir_weight[167][49],
reservoir_weight[167][50],
reservoir_weight[167][51],
reservoir_weight[167][52],
reservoir_weight[167][53],
reservoir_weight[167][54],
reservoir_weight[167][55],
reservoir_weight[167][56],
reservoir_weight[167][57],
reservoir_weight[167][58],
reservoir_weight[167][59],
reservoir_weight[167][60],
reservoir_weight[167][61],
reservoir_weight[167][62],
reservoir_weight[167][63],
reservoir_weight[167][64],
reservoir_weight[167][65],
reservoir_weight[167][66],
reservoir_weight[167][67],
reservoir_weight[167][68],
reservoir_weight[167][69],
reservoir_weight[167][70],
reservoir_weight[167][71],
reservoir_weight[167][72],
reservoir_weight[167][73],
reservoir_weight[167][74],
reservoir_weight[167][75],
reservoir_weight[167][76],
reservoir_weight[167][77],
reservoir_weight[167][78],
reservoir_weight[167][79],
reservoir_weight[167][80],
reservoir_weight[167][81],
reservoir_weight[167][82],
reservoir_weight[167][83],
reservoir_weight[167][84],
reservoir_weight[167][85],
reservoir_weight[167][86],
reservoir_weight[167][87],
reservoir_weight[167][88],
reservoir_weight[167][89],
reservoir_weight[167][90],
reservoir_weight[167][91],
reservoir_weight[167][92],
reservoir_weight[167][93],
reservoir_weight[167][94],
reservoir_weight[167][95],
reservoir_weight[167][96],
reservoir_weight[167][97],
reservoir_weight[167][98],
reservoir_weight[167][99],
reservoir_weight[167][100],
reservoir_weight[167][101],
reservoir_weight[167][102],
reservoir_weight[167][103],
reservoir_weight[167][104],
reservoir_weight[167][105],
reservoir_weight[167][106],
reservoir_weight[167][107],
reservoir_weight[167][108],
reservoir_weight[167][109],
reservoir_weight[167][110],
reservoir_weight[167][111],
reservoir_weight[167][112],
reservoir_weight[167][113],
reservoir_weight[167][114],
reservoir_weight[167][115],
reservoir_weight[167][116],
reservoir_weight[167][117],
reservoir_weight[167][118],
reservoir_weight[167][119],
reservoir_weight[167][120],
reservoir_weight[167][121],
reservoir_weight[167][122],
reservoir_weight[167][123],
reservoir_weight[167][124],
reservoir_weight[167][125],
reservoir_weight[167][126],
reservoir_weight[167][127],
reservoir_weight[167][128],
reservoir_weight[167][129],
reservoir_weight[167][130],
reservoir_weight[167][131],
reservoir_weight[167][132],
reservoir_weight[167][133],
reservoir_weight[167][134],
reservoir_weight[167][135],
reservoir_weight[167][136],
reservoir_weight[167][137],
reservoir_weight[167][138],
reservoir_weight[167][139],
reservoir_weight[167][140],
reservoir_weight[167][141],
reservoir_weight[167][142],
reservoir_weight[167][143],
reservoir_weight[167][144],
reservoir_weight[167][145],
reservoir_weight[167][146],
reservoir_weight[167][147],
reservoir_weight[167][148],
reservoir_weight[167][149],
reservoir_weight[167][150],
reservoir_weight[167][151],
reservoir_weight[167][152],
reservoir_weight[167][153],
reservoir_weight[167][154],
reservoir_weight[167][155],
reservoir_weight[167][156],
reservoir_weight[167][157],
reservoir_weight[167][158],
reservoir_weight[167][159],
reservoir_weight[167][160],
reservoir_weight[167][161],
reservoir_weight[167][162],
reservoir_weight[167][163],
reservoir_weight[167][164],
reservoir_weight[167][165],
reservoir_weight[167][166],
reservoir_weight[167][167],
reservoir_weight[167][168],
reservoir_weight[167][169],
reservoir_weight[167][170],
reservoir_weight[167][171],
reservoir_weight[167][172],
reservoir_weight[167][173],
reservoir_weight[167][174],
reservoir_weight[167][175],
reservoir_weight[167][176],
reservoir_weight[167][177],
reservoir_weight[167][178],
reservoir_weight[167][179],
reservoir_weight[167][180],
reservoir_weight[167][181],
reservoir_weight[167][182],
reservoir_weight[167][183],
reservoir_weight[167][184],
reservoir_weight[167][185],
reservoir_weight[167][186],
reservoir_weight[167][187],
reservoir_weight[167][188],
reservoir_weight[167][189],
reservoir_weight[167][190],
reservoir_weight[167][191],
reservoir_weight[167][192],
reservoir_weight[167][193],
reservoir_weight[167][194],
reservoir_weight[167][195],
reservoir_weight[167][196],
reservoir_weight[167][197],
reservoir_weight[167][198],
reservoir_weight[167][199]
},
{reservoir_weight[168][0],
reservoir_weight[168][1],
reservoir_weight[168][2],
reservoir_weight[168][3],
reservoir_weight[168][4],
reservoir_weight[168][5],
reservoir_weight[168][6],
reservoir_weight[168][7],
reservoir_weight[168][8],
reservoir_weight[168][9],
reservoir_weight[168][10],
reservoir_weight[168][11],
reservoir_weight[168][12],
reservoir_weight[168][13],
reservoir_weight[168][14],
reservoir_weight[168][15],
reservoir_weight[168][16],
reservoir_weight[168][17],
reservoir_weight[168][18],
reservoir_weight[168][19],
reservoir_weight[168][20],
reservoir_weight[168][21],
reservoir_weight[168][22],
reservoir_weight[168][23],
reservoir_weight[168][24],
reservoir_weight[168][25],
reservoir_weight[168][26],
reservoir_weight[168][27],
reservoir_weight[168][28],
reservoir_weight[168][29],
reservoir_weight[168][30],
reservoir_weight[168][31],
reservoir_weight[168][32],
reservoir_weight[168][33],
reservoir_weight[168][34],
reservoir_weight[168][35],
reservoir_weight[168][36],
reservoir_weight[168][37],
reservoir_weight[168][38],
reservoir_weight[168][39],
reservoir_weight[168][40],
reservoir_weight[168][41],
reservoir_weight[168][42],
reservoir_weight[168][43],
reservoir_weight[168][44],
reservoir_weight[168][45],
reservoir_weight[168][46],
reservoir_weight[168][47],
reservoir_weight[168][48],
reservoir_weight[168][49],
reservoir_weight[168][50],
reservoir_weight[168][51],
reservoir_weight[168][52],
reservoir_weight[168][53],
reservoir_weight[168][54],
reservoir_weight[168][55],
reservoir_weight[168][56],
reservoir_weight[168][57],
reservoir_weight[168][58],
reservoir_weight[168][59],
reservoir_weight[168][60],
reservoir_weight[168][61],
reservoir_weight[168][62],
reservoir_weight[168][63],
reservoir_weight[168][64],
reservoir_weight[168][65],
reservoir_weight[168][66],
reservoir_weight[168][67],
reservoir_weight[168][68],
reservoir_weight[168][69],
reservoir_weight[168][70],
reservoir_weight[168][71],
reservoir_weight[168][72],
reservoir_weight[168][73],
reservoir_weight[168][74],
reservoir_weight[168][75],
reservoir_weight[168][76],
reservoir_weight[168][77],
reservoir_weight[168][78],
reservoir_weight[168][79],
reservoir_weight[168][80],
reservoir_weight[168][81],
reservoir_weight[168][82],
reservoir_weight[168][83],
reservoir_weight[168][84],
reservoir_weight[168][85],
reservoir_weight[168][86],
reservoir_weight[168][87],
reservoir_weight[168][88],
reservoir_weight[168][89],
reservoir_weight[168][90],
reservoir_weight[168][91],
reservoir_weight[168][92],
reservoir_weight[168][93],
reservoir_weight[168][94],
reservoir_weight[168][95],
reservoir_weight[168][96],
reservoir_weight[168][97],
reservoir_weight[168][98],
reservoir_weight[168][99],
reservoir_weight[168][100],
reservoir_weight[168][101],
reservoir_weight[168][102],
reservoir_weight[168][103],
reservoir_weight[168][104],
reservoir_weight[168][105],
reservoir_weight[168][106],
reservoir_weight[168][107],
reservoir_weight[168][108],
reservoir_weight[168][109],
reservoir_weight[168][110],
reservoir_weight[168][111],
reservoir_weight[168][112],
reservoir_weight[168][113],
reservoir_weight[168][114],
reservoir_weight[168][115],
reservoir_weight[168][116],
reservoir_weight[168][117],
reservoir_weight[168][118],
reservoir_weight[168][119],
reservoir_weight[168][120],
reservoir_weight[168][121],
reservoir_weight[168][122],
reservoir_weight[168][123],
reservoir_weight[168][124],
reservoir_weight[168][125],
reservoir_weight[168][126],
reservoir_weight[168][127],
reservoir_weight[168][128],
reservoir_weight[168][129],
reservoir_weight[168][130],
reservoir_weight[168][131],
reservoir_weight[168][132],
reservoir_weight[168][133],
reservoir_weight[168][134],
reservoir_weight[168][135],
reservoir_weight[168][136],
reservoir_weight[168][137],
reservoir_weight[168][138],
reservoir_weight[168][139],
reservoir_weight[168][140],
reservoir_weight[168][141],
reservoir_weight[168][142],
reservoir_weight[168][143],
reservoir_weight[168][144],
reservoir_weight[168][145],
reservoir_weight[168][146],
reservoir_weight[168][147],
reservoir_weight[168][148],
reservoir_weight[168][149],
reservoir_weight[168][150],
reservoir_weight[168][151],
reservoir_weight[168][152],
reservoir_weight[168][153],
reservoir_weight[168][154],
reservoir_weight[168][155],
reservoir_weight[168][156],
reservoir_weight[168][157],
reservoir_weight[168][158],
reservoir_weight[168][159],
reservoir_weight[168][160],
reservoir_weight[168][161],
reservoir_weight[168][162],
reservoir_weight[168][163],
reservoir_weight[168][164],
reservoir_weight[168][165],
reservoir_weight[168][166],
reservoir_weight[168][167],
reservoir_weight[168][168],
reservoir_weight[168][169],
reservoir_weight[168][170],
reservoir_weight[168][171],
reservoir_weight[168][172],
reservoir_weight[168][173],
reservoir_weight[168][174],
reservoir_weight[168][175],
reservoir_weight[168][176],
reservoir_weight[168][177],
reservoir_weight[168][178],
reservoir_weight[168][179],
reservoir_weight[168][180],
reservoir_weight[168][181],
reservoir_weight[168][182],
reservoir_weight[168][183],
reservoir_weight[168][184],
reservoir_weight[168][185],
reservoir_weight[168][186],
reservoir_weight[168][187],
reservoir_weight[168][188],
reservoir_weight[168][189],
reservoir_weight[168][190],
reservoir_weight[168][191],
reservoir_weight[168][192],
reservoir_weight[168][193],
reservoir_weight[168][194],
reservoir_weight[168][195],
reservoir_weight[168][196],
reservoir_weight[168][197],
reservoir_weight[168][198],
reservoir_weight[168][199]
},
{reservoir_weight[169][0],
reservoir_weight[169][1],
reservoir_weight[169][2],
reservoir_weight[169][3],
reservoir_weight[169][4],
reservoir_weight[169][5],
reservoir_weight[169][6],
reservoir_weight[169][7],
reservoir_weight[169][8],
reservoir_weight[169][9],
reservoir_weight[169][10],
reservoir_weight[169][11],
reservoir_weight[169][12],
reservoir_weight[169][13],
reservoir_weight[169][14],
reservoir_weight[169][15],
reservoir_weight[169][16],
reservoir_weight[169][17],
reservoir_weight[169][18],
reservoir_weight[169][19],
reservoir_weight[169][20],
reservoir_weight[169][21],
reservoir_weight[169][22],
reservoir_weight[169][23],
reservoir_weight[169][24],
reservoir_weight[169][25],
reservoir_weight[169][26],
reservoir_weight[169][27],
reservoir_weight[169][28],
reservoir_weight[169][29],
reservoir_weight[169][30],
reservoir_weight[169][31],
reservoir_weight[169][32],
reservoir_weight[169][33],
reservoir_weight[169][34],
reservoir_weight[169][35],
reservoir_weight[169][36],
reservoir_weight[169][37],
reservoir_weight[169][38],
reservoir_weight[169][39],
reservoir_weight[169][40],
reservoir_weight[169][41],
reservoir_weight[169][42],
reservoir_weight[169][43],
reservoir_weight[169][44],
reservoir_weight[169][45],
reservoir_weight[169][46],
reservoir_weight[169][47],
reservoir_weight[169][48],
reservoir_weight[169][49],
reservoir_weight[169][50],
reservoir_weight[169][51],
reservoir_weight[169][52],
reservoir_weight[169][53],
reservoir_weight[169][54],
reservoir_weight[169][55],
reservoir_weight[169][56],
reservoir_weight[169][57],
reservoir_weight[169][58],
reservoir_weight[169][59],
reservoir_weight[169][60],
reservoir_weight[169][61],
reservoir_weight[169][62],
reservoir_weight[169][63],
reservoir_weight[169][64],
reservoir_weight[169][65],
reservoir_weight[169][66],
reservoir_weight[169][67],
reservoir_weight[169][68],
reservoir_weight[169][69],
reservoir_weight[169][70],
reservoir_weight[169][71],
reservoir_weight[169][72],
reservoir_weight[169][73],
reservoir_weight[169][74],
reservoir_weight[169][75],
reservoir_weight[169][76],
reservoir_weight[169][77],
reservoir_weight[169][78],
reservoir_weight[169][79],
reservoir_weight[169][80],
reservoir_weight[169][81],
reservoir_weight[169][82],
reservoir_weight[169][83],
reservoir_weight[169][84],
reservoir_weight[169][85],
reservoir_weight[169][86],
reservoir_weight[169][87],
reservoir_weight[169][88],
reservoir_weight[169][89],
reservoir_weight[169][90],
reservoir_weight[169][91],
reservoir_weight[169][92],
reservoir_weight[169][93],
reservoir_weight[169][94],
reservoir_weight[169][95],
reservoir_weight[169][96],
reservoir_weight[169][97],
reservoir_weight[169][98],
reservoir_weight[169][99],
reservoir_weight[169][100],
reservoir_weight[169][101],
reservoir_weight[169][102],
reservoir_weight[169][103],
reservoir_weight[169][104],
reservoir_weight[169][105],
reservoir_weight[169][106],
reservoir_weight[169][107],
reservoir_weight[169][108],
reservoir_weight[169][109],
reservoir_weight[169][110],
reservoir_weight[169][111],
reservoir_weight[169][112],
reservoir_weight[169][113],
reservoir_weight[169][114],
reservoir_weight[169][115],
reservoir_weight[169][116],
reservoir_weight[169][117],
reservoir_weight[169][118],
reservoir_weight[169][119],
reservoir_weight[169][120],
reservoir_weight[169][121],
reservoir_weight[169][122],
reservoir_weight[169][123],
reservoir_weight[169][124],
reservoir_weight[169][125],
reservoir_weight[169][126],
reservoir_weight[169][127],
reservoir_weight[169][128],
reservoir_weight[169][129],
reservoir_weight[169][130],
reservoir_weight[169][131],
reservoir_weight[169][132],
reservoir_weight[169][133],
reservoir_weight[169][134],
reservoir_weight[169][135],
reservoir_weight[169][136],
reservoir_weight[169][137],
reservoir_weight[169][138],
reservoir_weight[169][139],
reservoir_weight[169][140],
reservoir_weight[169][141],
reservoir_weight[169][142],
reservoir_weight[169][143],
reservoir_weight[169][144],
reservoir_weight[169][145],
reservoir_weight[169][146],
reservoir_weight[169][147],
reservoir_weight[169][148],
reservoir_weight[169][149],
reservoir_weight[169][150],
reservoir_weight[169][151],
reservoir_weight[169][152],
reservoir_weight[169][153],
reservoir_weight[169][154],
reservoir_weight[169][155],
reservoir_weight[169][156],
reservoir_weight[169][157],
reservoir_weight[169][158],
reservoir_weight[169][159],
reservoir_weight[169][160],
reservoir_weight[169][161],
reservoir_weight[169][162],
reservoir_weight[169][163],
reservoir_weight[169][164],
reservoir_weight[169][165],
reservoir_weight[169][166],
reservoir_weight[169][167],
reservoir_weight[169][168],
reservoir_weight[169][169],
reservoir_weight[169][170],
reservoir_weight[169][171],
reservoir_weight[169][172],
reservoir_weight[169][173],
reservoir_weight[169][174],
reservoir_weight[169][175],
reservoir_weight[169][176],
reservoir_weight[169][177],
reservoir_weight[169][178],
reservoir_weight[169][179],
reservoir_weight[169][180],
reservoir_weight[169][181],
reservoir_weight[169][182],
reservoir_weight[169][183],
reservoir_weight[169][184],
reservoir_weight[169][185],
reservoir_weight[169][186],
reservoir_weight[169][187],
reservoir_weight[169][188],
reservoir_weight[169][189],
reservoir_weight[169][190],
reservoir_weight[169][191],
reservoir_weight[169][192],
reservoir_weight[169][193],
reservoir_weight[169][194],
reservoir_weight[169][195],
reservoir_weight[169][196],
reservoir_weight[169][197],
reservoir_weight[169][198],
reservoir_weight[169][199]
},
{reservoir_weight[170][0],
reservoir_weight[170][1],
reservoir_weight[170][2],
reservoir_weight[170][3],
reservoir_weight[170][4],
reservoir_weight[170][5],
reservoir_weight[170][6],
reservoir_weight[170][7],
reservoir_weight[170][8],
reservoir_weight[170][9],
reservoir_weight[170][10],
reservoir_weight[170][11],
reservoir_weight[170][12],
reservoir_weight[170][13],
reservoir_weight[170][14],
reservoir_weight[170][15],
reservoir_weight[170][16],
reservoir_weight[170][17],
reservoir_weight[170][18],
reservoir_weight[170][19],
reservoir_weight[170][20],
reservoir_weight[170][21],
reservoir_weight[170][22],
reservoir_weight[170][23],
reservoir_weight[170][24],
reservoir_weight[170][25],
reservoir_weight[170][26],
reservoir_weight[170][27],
reservoir_weight[170][28],
reservoir_weight[170][29],
reservoir_weight[170][30],
reservoir_weight[170][31],
reservoir_weight[170][32],
reservoir_weight[170][33],
reservoir_weight[170][34],
reservoir_weight[170][35],
reservoir_weight[170][36],
reservoir_weight[170][37],
reservoir_weight[170][38],
reservoir_weight[170][39],
reservoir_weight[170][40],
reservoir_weight[170][41],
reservoir_weight[170][42],
reservoir_weight[170][43],
reservoir_weight[170][44],
reservoir_weight[170][45],
reservoir_weight[170][46],
reservoir_weight[170][47],
reservoir_weight[170][48],
reservoir_weight[170][49],
reservoir_weight[170][50],
reservoir_weight[170][51],
reservoir_weight[170][52],
reservoir_weight[170][53],
reservoir_weight[170][54],
reservoir_weight[170][55],
reservoir_weight[170][56],
reservoir_weight[170][57],
reservoir_weight[170][58],
reservoir_weight[170][59],
reservoir_weight[170][60],
reservoir_weight[170][61],
reservoir_weight[170][62],
reservoir_weight[170][63],
reservoir_weight[170][64],
reservoir_weight[170][65],
reservoir_weight[170][66],
reservoir_weight[170][67],
reservoir_weight[170][68],
reservoir_weight[170][69],
reservoir_weight[170][70],
reservoir_weight[170][71],
reservoir_weight[170][72],
reservoir_weight[170][73],
reservoir_weight[170][74],
reservoir_weight[170][75],
reservoir_weight[170][76],
reservoir_weight[170][77],
reservoir_weight[170][78],
reservoir_weight[170][79],
reservoir_weight[170][80],
reservoir_weight[170][81],
reservoir_weight[170][82],
reservoir_weight[170][83],
reservoir_weight[170][84],
reservoir_weight[170][85],
reservoir_weight[170][86],
reservoir_weight[170][87],
reservoir_weight[170][88],
reservoir_weight[170][89],
reservoir_weight[170][90],
reservoir_weight[170][91],
reservoir_weight[170][92],
reservoir_weight[170][93],
reservoir_weight[170][94],
reservoir_weight[170][95],
reservoir_weight[170][96],
reservoir_weight[170][97],
reservoir_weight[170][98],
reservoir_weight[170][99],
reservoir_weight[170][100],
reservoir_weight[170][101],
reservoir_weight[170][102],
reservoir_weight[170][103],
reservoir_weight[170][104],
reservoir_weight[170][105],
reservoir_weight[170][106],
reservoir_weight[170][107],
reservoir_weight[170][108],
reservoir_weight[170][109],
reservoir_weight[170][110],
reservoir_weight[170][111],
reservoir_weight[170][112],
reservoir_weight[170][113],
reservoir_weight[170][114],
reservoir_weight[170][115],
reservoir_weight[170][116],
reservoir_weight[170][117],
reservoir_weight[170][118],
reservoir_weight[170][119],
reservoir_weight[170][120],
reservoir_weight[170][121],
reservoir_weight[170][122],
reservoir_weight[170][123],
reservoir_weight[170][124],
reservoir_weight[170][125],
reservoir_weight[170][126],
reservoir_weight[170][127],
reservoir_weight[170][128],
reservoir_weight[170][129],
reservoir_weight[170][130],
reservoir_weight[170][131],
reservoir_weight[170][132],
reservoir_weight[170][133],
reservoir_weight[170][134],
reservoir_weight[170][135],
reservoir_weight[170][136],
reservoir_weight[170][137],
reservoir_weight[170][138],
reservoir_weight[170][139],
reservoir_weight[170][140],
reservoir_weight[170][141],
reservoir_weight[170][142],
reservoir_weight[170][143],
reservoir_weight[170][144],
reservoir_weight[170][145],
reservoir_weight[170][146],
reservoir_weight[170][147],
reservoir_weight[170][148],
reservoir_weight[170][149],
reservoir_weight[170][150],
reservoir_weight[170][151],
reservoir_weight[170][152],
reservoir_weight[170][153],
reservoir_weight[170][154],
reservoir_weight[170][155],
reservoir_weight[170][156],
reservoir_weight[170][157],
reservoir_weight[170][158],
reservoir_weight[170][159],
reservoir_weight[170][160],
reservoir_weight[170][161],
reservoir_weight[170][162],
reservoir_weight[170][163],
reservoir_weight[170][164],
reservoir_weight[170][165],
reservoir_weight[170][166],
reservoir_weight[170][167],
reservoir_weight[170][168],
reservoir_weight[170][169],
reservoir_weight[170][170],
reservoir_weight[170][171],
reservoir_weight[170][172],
reservoir_weight[170][173],
reservoir_weight[170][174],
reservoir_weight[170][175],
reservoir_weight[170][176],
reservoir_weight[170][177],
reservoir_weight[170][178],
reservoir_weight[170][179],
reservoir_weight[170][180],
reservoir_weight[170][181],
reservoir_weight[170][182],
reservoir_weight[170][183],
reservoir_weight[170][184],
reservoir_weight[170][185],
reservoir_weight[170][186],
reservoir_weight[170][187],
reservoir_weight[170][188],
reservoir_weight[170][189],
reservoir_weight[170][190],
reservoir_weight[170][191],
reservoir_weight[170][192],
reservoir_weight[170][193],
reservoir_weight[170][194],
reservoir_weight[170][195],
reservoir_weight[170][196],
reservoir_weight[170][197],
reservoir_weight[170][198],
reservoir_weight[170][199]
},
{reservoir_weight[171][0],
reservoir_weight[171][1],
reservoir_weight[171][2],
reservoir_weight[171][3],
reservoir_weight[171][4],
reservoir_weight[171][5],
reservoir_weight[171][6],
reservoir_weight[171][7],
reservoir_weight[171][8],
reservoir_weight[171][9],
reservoir_weight[171][10],
reservoir_weight[171][11],
reservoir_weight[171][12],
reservoir_weight[171][13],
reservoir_weight[171][14],
reservoir_weight[171][15],
reservoir_weight[171][16],
reservoir_weight[171][17],
reservoir_weight[171][18],
reservoir_weight[171][19],
reservoir_weight[171][20],
reservoir_weight[171][21],
reservoir_weight[171][22],
reservoir_weight[171][23],
reservoir_weight[171][24],
reservoir_weight[171][25],
reservoir_weight[171][26],
reservoir_weight[171][27],
reservoir_weight[171][28],
reservoir_weight[171][29],
reservoir_weight[171][30],
reservoir_weight[171][31],
reservoir_weight[171][32],
reservoir_weight[171][33],
reservoir_weight[171][34],
reservoir_weight[171][35],
reservoir_weight[171][36],
reservoir_weight[171][37],
reservoir_weight[171][38],
reservoir_weight[171][39],
reservoir_weight[171][40],
reservoir_weight[171][41],
reservoir_weight[171][42],
reservoir_weight[171][43],
reservoir_weight[171][44],
reservoir_weight[171][45],
reservoir_weight[171][46],
reservoir_weight[171][47],
reservoir_weight[171][48],
reservoir_weight[171][49],
reservoir_weight[171][50],
reservoir_weight[171][51],
reservoir_weight[171][52],
reservoir_weight[171][53],
reservoir_weight[171][54],
reservoir_weight[171][55],
reservoir_weight[171][56],
reservoir_weight[171][57],
reservoir_weight[171][58],
reservoir_weight[171][59],
reservoir_weight[171][60],
reservoir_weight[171][61],
reservoir_weight[171][62],
reservoir_weight[171][63],
reservoir_weight[171][64],
reservoir_weight[171][65],
reservoir_weight[171][66],
reservoir_weight[171][67],
reservoir_weight[171][68],
reservoir_weight[171][69],
reservoir_weight[171][70],
reservoir_weight[171][71],
reservoir_weight[171][72],
reservoir_weight[171][73],
reservoir_weight[171][74],
reservoir_weight[171][75],
reservoir_weight[171][76],
reservoir_weight[171][77],
reservoir_weight[171][78],
reservoir_weight[171][79],
reservoir_weight[171][80],
reservoir_weight[171][81],
reservoir_weight[171][82],
reservoir_weight[171][83],
reservoir_weight[171][84],
reservoir_weight[171][85],
reservoir_weight[171][86],
reservoir_weight[171][87],
reservoir_weight[171][88],
reservoir_weight[171][89],
reservoir_weight[171][90],
reservoir_weight[171][91],
reservoir_weight[171][92],
reservoir_weight[171][93],
reservoir_weight[171][94],
reservoir_weight[171][95],
reservoir_weight[171][96],
reservoir_weight[171][97],
reservoir_weight[171][98],
reservoir_weight[171][99],
reservoir_weight[171][100],
reservoir_weight[171][101],
reservoir_weight[171][102],
reservoir_weight[171][103],
reservoir_weight[171][104],
reservoir_weight[171][105],
reservoir_weight[171][106],
reservoir_weight[171][107],
reservoir_weight[171][108],
reservoir_weight[171][109],
reservoir_weight[171][110],
reservoir_weight[171][111],
reservoir_weight[171][112],
reservoir_weight[171][113],
reservoir_weight[171][114],
reservoir_weight[171][115],
reservoir_weight[171][116],
reservoir_weight[171][117],
reservoir_weight[171][118],
reservoir_weight[171][119],
reservoir_weight[171][120],
reservoir_weight[171][121],
reservoir_weight[171][122],
reservoir_weight[171][123],
reservoir_weight[171][124],
reservoir_weight[171][125],
reservoir_weight[171][126],
reservoir_weight[171][127],
reservoir_weight[171][128],
reservoir_weight[171][129],
reservoir_weight[171][130],
reservoir_weight[171][131],
reservoir_weight[171][132],
reservoir_weight[171][133],
reservoir_weight[171][134],
reservoir_weight[171][135],
reservoir_weight[171][136],
reservoir_weight[171][137],
reservoir_weight[171][138],
reservoir_weight[171][139],
reservoir_weight[171][140],
reservoir_weight[171][141],
reservoir_weight[171][142],
reservoir_weight[171][143],
reservoir_weight[171][144],
reservoir_weight[171][145],
reservoir_weight[171][146],
reservoir_weight[171][147],
reservoir_weight[171][148],
reservoir_weight[171][149],
reservoir_weight[171][150],
reservoir_weight[171][151],
reservoir_weight[171][152],
reservoir_weight[171][153],
reservoir_weight[171][154],
reservoir_weight[171][155],
reservoir_weight[171][156],
reservoir_weight[171][157],
reservoir_weight[171][158],
reservoir_weight[171][159],
reservoir_weight[171][160],
reservoir_weight[171][161],
reservoir_weight[171][162],
reservoir_weight[171][163],
reservoir_weight[171][164],
reservoir_weight[171][165],
reservoir_weight[171][166],
reservoir_weight[171][167],
reservoir_weight[171][168],
reservoir_weight[171][169],
reservoir_weight[171][170],
reservoir_weight[171][171],
reservoir_weight[171][172],
reservoir_weight[171][173],
reservoir_weight[171][174],
reservoir_weight[171][175],
reservoir_weight[171][176],
reservoir_weight[171][177],
reservoir_weight[171][178],
reservoir_weight[171][179],
reservoir_weight[171][180],
reservoir_weight[171][181],
reservoir_weight[171][182],
reservoir_weight[171][183],
reservoir_weight[171][184],
reservoir_weight[171][185],
reservoir_weight[171][186],
reservoir_weight[171][187],
reservoir_weight[171][188],
reservoir_weight[171][189],
reservoir_weight[171][190],
reservoir_weight[171][191],
reservoir_weight[171][192],
reservoir_weight[171][193],
reservoir_weight[171][194],
reservoir_weight[171][195],
reservoir_weight[171][196],
reservoir_weight[171][197],
reservoir_weight[171][198],
reservoir_weight[171][199]
},
{reservoir_weight[172][0],
reservoir_weight[172][1],
reservoir_weight[172][2],
reservoir_weight[172][3],
reservoir_weight[172][4],
reservoir_weight[172][5],
reservoir_weight[172][6],
reservoir_weight[172][7],
reservoir_weight[172][8],
reservoir_weight[172][9],
reservoir_weight[172][10],
reservoir_weight[172][11],
reservoir_weight[172][12],
reservoir_weight[172][13],
reservoir_weight[172][14],
reservoir_weight[172][15],
reservoir_weight[172][16],
reservoir_weight[172][17],
reservoir_weight[172][18],
reservoir_weight[172][19],
reservoir_weight[172][20],
reservoir_weight[172][21],
reservoir_weight[172][22],
reservoir_weight[172][23],
reservoir_weight[172][24],
reservoir_weight[172][25],
reservoir_weight[172][26],
reservoir_weight[172][27],
reservoir_weight[172][28],
reservoir_weight[172][29],
reservoir_weight[172][30],
reservoir_weight[172][31],
reservoir_weight[172][32],
reservoir_weight[172][33],
reservoir_weight[172][34],
reservoir_weight[172][35],
reservoir_weight[172][36],
reservoir_weight[172][37],
reservoir_weight[172][38],
reservoir_weight[172][39],
reservoir_weight[172][40],
reservoir_weight[172][41],
reservoir_weight[172][42],
reservoir_weight[172][43],
reservoir_weight[172][44],
reservoir_weight[172][45],
reservoir_weight[172][46],
reservoir_weight[172][47],
reservoir_weight[172][48],
reservoir_weight[172][49],
reservoir_weight[172][50],
reservoir_weight[172][51],
reservoir_weight[172][52],
reservoir_weight[172][53],
reservoir_weight[172][54],
reservoir_weight[172][55],
reservoir_weight[172][56],
reservoir_weight[172][57],
reservoir_weight[172][58],
reservoir_weight[172][59],
reservoir_weight[172][60],
reservoir_weight[172][61],
reservoir_weight[172][62],
reservoir_weight[172][63],
reservoir_weight[172][64],
reservoir_weight[172][65],
reservoir_weight[172][66],
reservoir_weight[172][67],
reservoir_weight[172][68],
reservoir_weight[172][69],
reservoir_weight[172][70],
reservoir_weight[172][71],
reservoir_weight[172][72],
reservoir_weight[172][73],
reservoir_weight[172][74],
reservoir_weight[172][75],
reservoir_weight[172][76],
reservoir_weight[172][77],
reservoir_weight[172][78],
reservoir_weight[172][79],
reservoir_weight[172][80],
reservoir_weight[172][81],
reservoir_weight[172][82],
reservoir_weight[172][83],
reservoir_weight[172][84],
reservoir_weight[172][85],
reservoir_weight[172][86],
reservoir_weight[172][87],
reservoir_weight[172][88],
reservoir_weight[172][89],
reservoir_weight[172][90],
reservoir_weight[172][91],
reservoir_weight[172][92],
reservoir_weight[172][93],
reservoir_weight[172][94],
reservoir_weight[172][95],
reservoir_weight[172][96],
reservoir_weight[172][97],
reservoir_weight[172][98],
reservoir_weight[172][99],
reservoir_weight[172][100],
reservoir_weight[172][101],
reservoir_weight[172][102],
reservoir_weight[172][103],
reservoir_weight[172][104],
reservoir_weight[172][105],
reservoir_weight[172][106],
reservoir_weight[172][107],
reservoir_weight[172][108],
reservoir_weight[172][109],
reservoir_weight[172][110],
reservoir_weight[172][111],
reservoir_weight[172][112],
reservoir_weight[172][113],
reservoir_weight[172][114],
reservoir_weight[172][115],
reservoir_weight[172][116],
reservoir_weight[172][117],
reservoir_weight[172][118],
reservoir_weight[172][119],
reservoir_weight[172][120],
reservoir_weight[172][121],
reservoir_weight[172][122],
reservoir_weight[172][123],
reservoir_weight[172][124],
reservoir_weight[172][125],
reservoir_weight[172][126],
reservoir_weight[172][127],
reservoir_weight[172][128],
reservoir_weight[172][129],
reservoir_weight[172][130],
reservoir_weight[172][131],
reservoir_weight[172][132],
reservoir_weight[172][133],
reservoir_weight[172][134],
reservoir_weight[172][135],
reservoir_weight[172][136],
reservoir_weight[172][137],
reservoir_weight[172][138],
reservoir_weight[172][139],
reservoir_weight[172][140],
reservoir_weight[172][141],
reservoir_weight[172][142],
reservoir_weight[172][143],
reservoir_weight[172][144],
reservoir_weight[172][145],
reservoir_weight[172][146],
reservoir_weight[172][147],
reservoir_weight[172][148],
reservoir_weight[172][149],
reservoir_weight[172][150],
reservoir_weight[172][151],
reservoir_weight[172][152],
reservoir_weight[172][153],
reservoir_weight[172][154],
reservoir_weight[172][155],
reservoir_weight[172][156],
reservoir_weight[172][157],
reservoir_weight[172][158],
reservoir_weight[172][159],
reservoir_weight[172][160],
reservoir_weight[172][161],
reservoir_weight[172][162],
reservoir_weight[172][163],
reservoir_weight[172][164],
reservoir_weight[172][165],
reservoir_weight[172][166],
reservoir_weight[172][167],
reservoir_weight[172][168],
reservoir_weight[172][169],
reservoir_weight[172][170],
reservoir_weight[172][171],
reservoir_weight[172][172],
reservoir_weight[172][173],
reservoir_weight[172][174],
reservoir_weight[172][175],
reservoir_weight[172][176],
reservoir_weight[172][177],
reservoir_weight[172][178],
reservoir_weight[172][179],
reservoir_weight[172][180],
reservoir_weight[172][181],
reservoir_weight[172][182],
reservoir_weight[172][183],
reservoir_weight[172][184],
reservoir_weight[172][185],
reservoir_weight[172][186],
reservoir_weight[172][187],
reservoir_weight[172][188],
reservoir_weight[172][189],
reservoir_weight[172][190],
reservoir_weight[172][191],
reservoir_weight[172][192],
reservoir_weight[172][193],
reservoir_weight[172][194],
reservoir_weight[172][195],
reservoir_weight[172][196],
reservoir_weight[172][197],
reservoir_weight[172][198],
reservoir_weight[172][199]
},
{reservoir_weight[173][0],
reservoir_weight[173][1],
reservoir_weight[173][2],
reservoir_weight[173][3],
reservoir_weight[173][4],
reservoir_weight[173][5],
reservoir_weight[173][6],
reservoir_weight[173][7],
reservoir_weight[173][8],
reservoir_weight[173][9],
reservoir_weight[173][10],
reservoir_weight[173][11],
reservoir_weight[173][12],
reservoir_weight[173][13],
reservoir_weight[173][14],
reservoir_weight[173][15],
reservoir_weight[173][16],
reservoir_weight[173][17],
reservoir_weight[173][18],
reservoir_weight[173][19],
reservoir_weight[173][20],
reservoir_weight[173][21],
reservoir_weight[173][22],
reservoir_weight[173][23],
reservoir_weight[173][24],
reservoir_weight[173][25],
reservoir_weight[173][26],
reservoir_weight[173][27],
reservoir_weight[173][28],
reservoir_weight[173][29],
reservoir_weight[173][30],
reservoir_weight[173][31],
reservoir_weight[173][32],
reservoir_weight[173][33],
reservoir_weight[173][34],
reservoir_weight[173][35],
reservoir_weight[173][36],
reservoir_weight[173][37],
reservoir_weight[173][38],
reservoir_weight[173][39],
reservoir_weight[173][40],
reservoir_weight[173][41],
reservoir_weight[173][42],
reservoir_weight[173][43],
reservoir_weight[173][44],
reservoir_weight[173][45],
reservoir_weight[173][46],
reservoir_weight[173][47],
reservoir_weight[173][48],
reservoir_weight[173][49],
reservoir_weight[173][50],
reservoir_weight[173][51],
reservoir_weight[173][52],
reservoir_weight[173][53],
reservoir_weight[173][54],
reservoir_weight[173][55],
reservoir_weight[173][56],
reservoir_weight[173][57],
reservoir_weight[173][58],
reservoir_weight[173][59],
reservoir_weight[173][60],
reservoir_weight[173][61],
reservoir_weight[173][62],
reservoir_weight[173][63],
reservoir_weight[173][64],
reservoir_weight[173][65],
reservoir_weight[173][66],
reservoir_weight[173][67],
reservoir_weight[173][68],
reservoir_weight[173][69],
reservoir_weight[173][70],
reservoir_weight[173][71],
reservoir_weight[173][72],
reservoir_weight[173][73],
reservoir_weight[173][74],
reservoir_weight[173][75],
reservoir_weight[173][76],
reservoir_weight[173][77],
reservoir_weight[173][78],
reservoir_weight[173][79],
reservoir_weight[173][80],
reservoir_weight[173][81],
reservoir_weight[173][82],
reservoir_weight[173][83],
reservoir_weight[173][84],
reservoir_weight[173][85],
reservoir_weight[173][86],
reservoir_weight[173][87],
reservoir_weight[173][88],
reservoir_weight[173][89],
reservoir_weight[173][90],
reservoir_weight[173][91],
reservoir_weight[173][92],
reservoir_weight[173][93],
reservoir_weight[173][94],
reservoir_weight[173][95],
reservoir_weight[173][96],
reservoir_weight[173][97],
reservoir_weight[173][98],
reservoir_weight[173][99],
reservoir_weight[173][100],
reservoir_weight[173][101],
reservoir_weight[173][102],
reservoir_weight[173][103],
reservoir_weight[173][104],
reservoir_weight[173][105],
reservoir_weight[173][106],
reservoir_weight[173][107],
reservoir_weight[173][108],
reservoir_weight[173][109],
reservoir_weight[173][110],
reservoir_weight[173][111],
reservoir_weight[173][112],
reservoir_weight[173][113],
reservoir_weight[173][114],
reservoir_weight[173][115],
reservoir_weight[173][116],
reservoir_weight[173][117],
reservoir_weight[173][118],
reservoir_weight[173][119],
reservoir_weight[173][120],
reservoir_weight[173][121],
reservoir_weight[173][122],
reservoir_weight[173][123],
reservoir_weight[173][124],
reservoir_weight[173][125],
reservoir_weight[173][126],
reservoir_weight[173][127],
reservoir_weight[173][128],
reservoir_weight[173][129],
reservoir_weight[173][130],
reservoir_weight[173][131],
reservoir_weight[173][132],
reservoir_weight[173][133],
reservoir_weight[173][134],
reservoir_weight[173][135],
reservoir_weight[173][136],
reservoir_weight[173][137],
reservoir_weight[173][138],
reservoir_weight[173][139],
reservoir_weight[173][140],
reservoir_weight[173][141],
reservoir_weight[173][142],
reservoir_weight[173][143],
reservoir_weight[173][144],
reservoir_weight[173][145],
reservoir_weight[173][146],
reservoir_weight[173][147],
reservoir_weight[173][148],
reservoir_weight[173][149],
reservoir_weight[173][150],
reservoir_weight[173][151],
reservoir_weight[173][152],
reservoir_weight[173][153],
reservoir_weight[173][154],
reservoir_weight[173][155],
reservoir_weight[173][156],
reservoir_weight[173][157],
reservoir_weight[173][158],
reservoir_weight[173][159],
reservoir_weight[173][160],
reservoir_weight[173][161],
reservoir_weight[173][162],
reservoir_weight[173][163],
reservoir_weight[173][164],
reservoir_weight[173][165],
reservoir_weight[173][166],
reservoir_weight[173][167],
reservoir_weight[173][168],
reservoir_weight[173][169],
reservoir_weight[173][170],
reservoir_weight[173][171],
reservoir_weight[173][172],
reservoir_weight[173][173],
reservoir_weight[173][174],
reservoir_weight[173][175],
reservoir_weight[173][176],
reservoir_weight[173][177],
reservoir_weight[173][178],
reservoir_weight[173][179],
reservoir_weight[173][180],
reservoir_weight[173][181],
reservoir_weight[173][182],
reservoir_weight[173][183],
reservoir_weight[173][184],
reservoir_weight[173][185],
reservoir_weight[173][186],
reservoir_weight[173][187],
reservoir_weight[173][188],
reservoir_weight[173][189],
reservoir_weight[173][190],
reservoir_weight[173][191],
reservoir_weight[173][192],
reservoir_weight[173][193],
reservoir_weight[173][194],
reservoir_weight[173][195],
reservoir_weight[173][196],
reservoir_weight[173][197],
reservoir_weight[173][198],
reservoir_weight[173][199]
},
{reservoir_weight[174][0],
reservoir_weight[174][1],
reservoir_weight[174][2],
reservoir_weight[174][3],
reservoir_weight[174][4],
reservoir_weight[174][5],
reservoir_weight[174][6],
reservoir_weight[174][7],
reservoir_weight[174][8],
reservoir_weight[174][9],
reservoir_weight[174][10],
reservoir_weight[174][11],
reservoir_weight[174][12],
reservoir_weight[174][13],
reservoir_weight[174][14],
reservoir_weight[174][15],
reservoir_weight[174][16],
reservoir_weight[174][17],
reservoir_weight[174][18],
reservoir_weight[174][19],
reservoir_weight[174][20],
reservoir_weight[174][21],
reservoir_weight[174][22],
reservoir_weight[174][23],
reservoir_weight[174][24],
reservoir_weight[174][25],
reservoir_weight[174][26],
reservoir_weight[174][27],
reservoir_weight[174][28],
reservoir_weight[174][29],
reservoir_weight[174][30],
reservoir_weight[174][31],
reservoir_weight[174][32],
reservoir_weight[174][33],
reservoir_weight[174][34],
reservoir_weight[174][35],
reservoir_weight[174][36],
reservoir_weight[174][37],
reservoir_weight[174][38],
reservoir_weight[174][39],
reservoir_weight[174][40],
reservoir_weight[174][41],
reservoir_weight[174][42],
reservoir_weight[174][43],
reservoir_weight[174][44],
reservoir_weight[174][45],
reservoir_weight[174][46],
reservoir_weight[174][47],
reservoir_weight[174][48],
reservoir_weight[174][49],
reservoir_weight[174][50],
reservoir_weight[174][51],
reservoir_weight[174][52],
reservoir_weight[174][53],
reservoir_weight[174][54],
reservoir_weight[174][55],
reservoir_weight[174][56],
reservoir_weight[174][57],
reservoir_weight[174][58],
reservoir_weight[174][59],
reservoir_weight[174][60],
reservoir_weight[174][61],
reservoir_weight[174][62],
reservoir_weight[174][63],
reservoir_weight[174][64],
reservoir_weight[174][65],
reservoir_weight[174][66],
reservoir_weight[174][67],
reservoir_weight[174][68],
reservoir_weight[174][69],
reservoir_weight[174][70],
reservoir_weight[174][71],
reservoir_weight[174][72],
reservoir_weight[174][73],
reservoir_weight[174][74],
reservoir_weight[174][75],
reservoir_weight[174][76],
reservoir_weight[174][77],
reservoir_weight[174][78],
reservoir_weight[174][79],
reservoir_weight[174][80],
reservoir_weight[174][81],
reservoir_weight[174][82],
reservoir_weight[174][83],
reservoir_weight[174][84],
reservoir_weight[174][85],
reservoir_weight[174][86],
reservoir_weight[174][87],
reservoir_weight[174][88],
reservoir_weight[174][89],
reservoir_weight[174][90],
reservoir_weight[174][91],
reservoir_weight[174][92],
reservoir_weight[174][93],
reservoir_weight[174][94],
reservoir_weight[174][95],
reservoir_weight[174][96],
reservoir_weight[174][97],
reservoir_weight[174][98],
reservoir_weight[174][99],
reservoir_weight[174][100],
reservoir_weight[174][101],
reservoir_weight[174][102],
reservoir_weight[174][103],
reservoir_weight[174][104],
reservoir_weight[174][105],
reservoir_weight[174][106],
reservoir_weight[174][107],
reservoir_weight[174][108],
reservoir_weight[174][109],
reservoir_weight[174][110],
reservoir_weight[174][111],
reservoir_weight[174][112],
reservoir_weight[174][113],
reservoir_weight[174][114],
reservoir_weight[174][115],
reservoir_weight[174][116],
reservoir_weight[174][117],
reservoir_weight[174][118],
reservoir_weight[174][119],
reservoir_weight[174][120],
reservoir_weight[174][121],
reservoir_weight[174][122],
reservoir_weight[174][123],
reservoir_weight[174][124],
reservoir_weight[174][125],
reservoir_weight[174][126],
reservoir_weight[174][127],
reservoir_weight[174][128],
reservoir_weight[174][129],
reservoir_weight[174][130],
reservoir_weight[174][131],
reservoir_weight[174][132],
reservoir_weight[174][133],
reservoir_weight[174][134],
reservoir_weight[174][135],
reservoir_weight[174][136],
reservoir_weight[174][137],
reservoir_weight[174][138],
reservoir_weight[174][139],
reservoir_weight[174][140],
reservoir_weight[174][141],
reservoir_weight[174][142],
reservoir_weight[174][143],
reservoir_weight[174][144],
reservoir_weight[174][145],
reservoir_weight[174][146],
reservoir_weight[174][147],
reservoir_weight[174][148],
reservoir_weight[174][149],
reservoir_weight[174][150],
reservoir_weight[174][151],
reservoir_weight[174][152],
reservoir_weight[174][153],
reservoir_weight[174][154],
reservoir_weight[174][155],
reservoir_weight[174][156],
reservoir_weight[174][157],
reservoir_weight[174][158],
reservoir_weight[174][159],
reservoir_weight[174][160],
reservoir_weight[174][161],
reservoir_weight[174][162],
reservoir_weight[174][163],
reservoir_weight[174][164],
reservoir_weight[174][165],
reservoir_weight[174][166],
reservoir_weight[174][167],
reservoir_weight[174][168],
reservoir_weight[174][169],
reservoir_weight[174][170],
reservoir_weight[174][171],
reservoir_weight[174][172],
reservoir_weight[174][173],
reservoir_weight[174][174],
reservoir_weight[174][175],
reservoir_weight[174][176],
reservoir_weight[174][177],
reservoir_weight[174][178],
reservoir_weight[174][179],
reservoir_weight[174][180],
reservoir_weight[174][181],
reservoir_weight[174][182],
reservoir_weight[174][183],
reservoir_weight[174][184],
reservoir_weight[174][185],
reservoir_weight[174][186],
reservoir_weight[174][187],
reservoir_weight[174][188],
reservoir_weight[174][189],
reservoir_weight[174][190],
reservoir_weight[174][191],
reservoir_weight[174][192],
reservoir_weight[174][193],
reservoir_weight[174][194],
reservoir_weight[174][195],
reservoir_weight[174][196],
reservoir_weight[174][197],
reservoir_weight[174][198],
reservoir_weight[174][199]
},
{reservoir_weight[175][0],
reservoir_weight[175][1],
reservoir_weight[175][2],
reservoir_weight[175][3],
reservoir_weight[175][4],
reservoir_weight[175][5],
reservoir_weight[175][6],
reservoir_weight[175][7],
reservoir_weight[175][8],
reservoir_weight[175][9],
reservoir_weight[175][10],
reservoir_weight[175][11],
reservoir_weight[175][12],
reservoir_weight[175][13],
reservoir_weight[175][14],
reservoir_weight[175][15],
reservoir_weight[175][16],
reservoir_weight[175][17],
reservoir_weight[175][18],
reservoir_weight[175][19],
reservoir_weight[175][20],
reservoir_weight[175][21],
reservoir_weight[175][22],
reservoir_weight[175][23],
reservoir_weight[175][24],
reservoir_weight[175][25],
reservoir_weight[175][26],
reservoir_weight[175][27],
reservoir_weight[175][28],
reservoir_weight[175][29],
reservoir_weight[175][30],
reservoir_weight[175][31],
reservoir_weight[175][32],
reservoir_weight[175][33],
reservoir_weight[175][34],
reservoir_weight[175][35],
reservoir_weight[175][36],
reservoir_weight[175][37],
reservoir_weight[175][38],
reservoir_weight[175][39],
reservoir_weight[175][40],
reservoir_weight[175][41],
reservoir_weight[175][42],
reservoir_weight[175][43],
reservoir_weight[175][44],
reservoir_weight[175][45],
reservoir_weight[175][46],
reservoir_weight[175][47],
reservoir_weight[175][48],
reservoir_weight[175][49],
reservoir_weight[175][50],
reservoir_weight[175][51],
reservoir_weight[175][52],
reservoir_weight[175][53],
reservoir_weight[175][54],
reservoir_weight[175][55],
reservoir_weight[175][56],
reservoir_weight[175][57],
reservoir_weight[175][58],
reservoir_weight[175][59],
reservoir_weight[175][60],
reservoir_weight[175][61],
reservoir_weight[175][62],
reservoir_weight[175][63],
reservoir_weight[175][64],
reservoir_weight[175][65],
reservoir_weight[175][66],
reservoir_weight[175][67],
reservoir_weight[175][68],
reservoir_weight[175][69],
reservoir_weight[175][70],
reservoir_weight[175][71],
reservoir_weight[175][72],
reservoir_weight[175][73],
reservoir_weight[175][74],
reservoir_weight[175][75],
reservoir_weight[175][76],
reservoir_weight[175][77],
reservoir_weight[175][78],
reservoir_weight[175][79],
reservoir_weight[175][80],
reservoir_weight[175][81],
reservoir_weight[175][82],
reservoir_weight[175][83],
reservoir_weight[175][84],
reservoir_weight[175][85],
reservoir_weight[175][86],
reservoir_weight[175][87],
reservoir_weight[175][88],
reservoir_weight[175][89],
reservoir_weight[175][90],
reservoir_weight[175][91],
reservoir_weight[175][92],
reservoir_weight[175][93],
reservoir_weight[175][94],
reservoir_weight[175][95],
reservoir_weight[175][96],
reservoir_weight[175][97],
reservoir_weight[175][98],
reservoir_weight[175][99],
reservoir_weight[175][100],
reservoir_weight[175][101],
reservoir_weight[175][102],
reservoir_weight[175][103],
reservoir_weight[175][104],
reservoir_weight[175][105],
reservoir_weight[175][106],
reservoir_weight[175][107],
reservoir_weight[175][108],
reservoir_weight[175][109],
reservoir_weight[175][110],
reservoir_weight[175][111],
reservoir_weight[175][112],
reservoir_weight[175][113],
reservoir_weight[175][114],
reservoir_weight[175][115],
reservoir_weight[175][116],
reservoir_weight[175][117],
reservoir_weight[175][118],
reservoir_weight[175][119],
reservoir_weight[175][120],
reservoir_weight[175][121],
reservoir_weight[175][122],
reservoir_weight[175][123],
reservoir_weight[175][124],
reservoir_weight[175][125],
reservoir_weight[175][126],
reservoir_weight[175][127],
reservoir_weight[175][128],
reservoir_weight[175][129],
reservoir_weight[175][130],
reservoir_weight[175][131],
reservoir_weight[175][132],
reservoir_weight[175][133],
reservoir_weight[175][134],
reservoir_weight[175][135],
reservoir_weight[175][136],
reservoir_weight[175][137],
reservoir_weight[175][138],
reservoir_weight[175][139],
reservoir_weight[175][140],
reservoir_weight[175][141],
reservoir_weight[175][142],
reservoir_weight[175][143],
reservoir_weight[175][144],
reservoir_weight[175][145],
reservoir_weight[175][146],
reservoir_weight[175][147],
reservoir_weight[175][148],
reservoir_weight[175][149],
reservoir_weight[175][150],
reservoir_weight[175][151],
reservoir_weight[175][152],
reservoir_weight[175][153],
reservoir_weight[175][154],
reservoir_weight[175][155],
reservoir_weight[175][156],
reservoir_weight[175][157],
reservoir_weight[175][158],
reservoir_weight[175][159],
reservoir_weight[175][160],
reservoir_weight[175][161],
reservoir_weight[175][162],
reservoir_weight[175][163],
reservoir_weight[175][164],
reservoir_weight[175][165],
reservoir_weight[175][166],
reservoir_weight[175][167],
reservoir_weight[175][168],
reservoir_weight[175][169],
reservoir_weight[175][170],
reservoir_weight[175][171],
reservoir_weight[175][172],
reservoir_weight[175][173],
reservoir_weight[175][174],
reservoir_weight[175][175],
reservoir_weight[175][176],
reservoir_weight[175][177],
reservoir_weight[175][178],
reservoir_weight[175][179],
reservoir_weight[175][180],
reservoir_weight[175][181],
reservoir_weight[175][182],
reservoir_weight[175][183],
reservoir_weight[175][184],
reservoir_weight[175][185],
reservoir_weight[175][186],
reservoir_weight[175][187],
reservoir_weight[175][188],
reservoir_weight[175][189],
reservoir_weight[175][190],
reservoir_weight[175][191],
reservoir_weight[175][192],
reservoir_weight[175][193],
reservoir_weight[175][194],
reservoir_weight[175][195],
reservoir_weight[175][196],
reservoir_weight[175][197],
reservoir_weight[175][198],
reservoir_weight[175][199]
},
{reservoir_weight[176][0],
reservoir_weight[176][1],
reservoir_weight[176][2],
reservoir_weight[176][3],
reservoir_weight[176][4],
reservoir_weight[176][5],
reservoir_weight[176][6],
reservoir_weight[176][7],
reservoir_weight[176][8],
reservoir_weight[176][9],
reservoir_weight[176][10],
reservoir_weight[176][11],
reservoir_weight[176][12],
reservoir_weight[176][13],
reservoir_weight[176][14],
reservoir_weight[176][15],
reservoir_weight[176][16],
reservoir_weight[176][17],
reservoir_weight[176][18],
reservoir_weight[176][19],
reservoir_weight[176][20],
reservoir_weight[176][21],
reservoir_weight[176][22],
reservoir_weight[176][23],
reservoir_weight[176][24],
reservoir_weight[176][25],
reservoir_weight[176][26],
reservoir_weight[176][27],
reservoir_weight[176][28],
reservoir_weight[176][29],
reservoir_weight[176][30],
reservoir_weight[176][31],
reservoir_weight[176][32],
reservoir_weight[176][33],
reservoir_weight[176][34],
reservoir_weight[176][35],
reservoir_weight[176][36],
reservoir_weight[176][37],
reservoir_weight[176][38],
reservoir_weight[176][39],
reservoir_weight[176][40],
reservoir_weight[176][41],
reservoir_weight[176][42],
reservoir_weight[176][43],
reservoir_weight[176][44],
reservoir_weight[176][45],
reservoir_weight[176][46],
reservoir_weight[176][47],
reservoir_weight[176][48],
reservoir_weight[176][49],
reservoir_weight[176][50],
reservoir_weight[176][51],
reservoir_weight[176][52],
reservoir_weight[176][53],
reservoir_weight[176][54],
reservoir_weight[176][55],
reservoir_weight[176][56],
reservoir_weight[176][57],
reservoir_weight[176][58],
reservoir_weight[176][59],
reservoir_weight[176][60],
reservoir_weight[176][61],
reservoir_weight[176][62],
reservoir_weight[176][63],
reservoir_weight[176][64],
reservoir_weight[176][65],
reservoir_weight[176][66],
reservoir_weight[176][67],
reservoir_weight[176][68],
reservoir_weight[176][69],
reservoir_weight[176][70],
reservoir_weight[176][71],
reservoir_weight[176][72],
reservoir_weight[176][73],
reservoir_weight[176][74],
reservoir_weight[176][75],
reservoir_weight[176][76],
reservoir_weight[176][77],
reservoir_weight[176][78],
reservoir_weight[176][79],
reservoir_weight[176][80],
reservoir_weight[176][81],
reservoir_weight[176][82],
reservoir_weight[176][83],
reservoir_weight[176][84],
reservoir_weight[176][85],
reservoir_weight[176][86],
reservoir_weight[176][87],
reservoir_weight[176][88],
reservoir_weight[176][89],
reservoir_weight[176][90],
reservoir_weight[176][91],
reservoir_weight[176][92],
reservoir_weight[176][93],
reservoir_weight[176][94],
reservoir_weight[176][95],
reservoir_weight[176][96],
reservoir_weight[176][97],
reservoir_weight[176][98],
reservoir_weight[176][99],
reservoir_weight[176][100],
reservoir_weight[176][101],
reservoir_weight[176][102],
reservoir_weight[176][103],
reservoir_weight[176][104],
reservoir_weight[176][105],
reservoir_weight[176][106],
reservoir_weight[176][107],
reservoir_weight[176][108],
reservoir_weight[176][109],
reservoir_weight[176][110],
reservoir_weight[176][111],
reservoir_weight[176][112],
reservoir_weight[176][113],
reservoir_weight[176][114],
reservoir_weight[176][115],
reservoir_weight[176][116],
reservoir_weight[176][117],
reservoir_weight[176][118],
reservoir_weight[176][119],
reservoir_weight[176][120],
reservoir_weight[176][121],
reservoir_weight[176][122],
reservoir_weight[176][123],
reservoir_weight[176][124],
reservoir_weight[176][125],
reservoir_weight[176][126],
reservoir_weight[176][127],
reservoir_weight[176][128],
reservoir_weight[176][129],
reservoir_weight[176][130],
reservoir_weight[176][131],
reservoir_weight[176][132],
reservoir_weight[176][133],
reservoir_weight[176][134],
reservoir_weight[176][135],
reservoir_weight[176][136],
reservoir_weight[176][137],
reservoir_weight[176][138],
reservoir_weight[176][139],
reservoir_weight[176][140],
reservoir_weight[176][141],
reservoir_weight[176][142],
reservoir_weight[176][143],
reservoir_weight[176][144],
reservoir_weight[176][145],
reservoir_weight[176][146],
reservoir_weight[176][147],
reservoir_weight[176][148],
reservoir_weight[176][149],
reservoir_weight[176][150],
reservoir_weight[176][151],
reservoir_weight[176][152],
reservoir_weight[176][153],
reservoir_weight[176][154],
reservoir_weight[176][155],
reservoir_weight[176][156],
reservoir_weight[176][157],
reservoir_weight[176][158],
reservoir_weight[176][159],
reservoir_weight[176][160],
reservoir_weight[176][161],
reservoir_weight[176][162],
reservoir_weight[176][163],
reservoir_weight[176][164],
reservoir_weight[176][165],
reservoir_weight[176][166],
reservoir_weight[176][167],
reservoir_weight[176][168],
reservoir_weight[176][169],
reservoir_weight[176][170],
reservoir_weight[176][171],
reservoir_weight[176][172],
reservoir_weight[176][173],
reservoir_weight[176][174],
reservoir_weight[176][175],
reservoir_weight[176][176],
reservoir_weight[176][177],
reservoir_weight[176][178],
reservoir_weight[176][179],
reservoir_weight[176][180],
reservoir_weight[176][181],
reservoir_weight[176][182],
reservoir_weight[176][183],
reservoir_weight[176][184],
reservoir_weight[176][185],
reservoir_weight[176][186],
reservoir_weight[176][187],
reservoir_weight[176][188],
reservoir_weight[176][189],
reservoir_weight[176][190],
reservoir_weight[176][191],
reservoir_weight[176][192],
reservoir_weight[176][193],
reservoir_weight[176][194],
reservoir_weight[176][195],
reservoir_weight[176][196],
reservoir_weight[176][197],
reservoir_weight[176][198],
reservoir_weight[176][199]
},
{reservoir_weight[177][0],
reservoir_weight[177][1],
reservoir_weight[177][2],
reservoir_weight[177][3],
reservoir_weight[177][4],
reservoir_weight[177][5],
reservoir_weight[177][6],
reservoir_weight[177][7],
reservoir_weight[177][8],
reservoir_weight[177][9],
reservoir_weight[177][10],
reservoir_weight[177][11],
reservoir_weight[177][12],
reservoir_weight[177][13],
reservoir_weight[177][14],
reservoir_weight[177][15],
reservoir_weight[177][16],
reservoir_weight[177][17],
reservoir_weight[177][18],
reservoir_weight[177][19],
reservoir_weight[177][20],
reservoir_weight[177][21],
reservoir_weight[177][22],
reservoir_weight[177][23],
reservoir_weight[177][24],
reservoir_weight[177][25],
reservoir_weight[177][26],
reservoir_weight[177][27],
reservoir_weight[177][28],
reservoir_weight[177][29],
reservoir_weight[177][30],
reservoir_weight[177][31],
reservoir_weight[177][32],
reservoir_weight[177][33],
reservoir_weight[177][34],
reservoir_weight[177][35],
reservoir_weight[177][36],
reservoir_weight[177][37],
reservoir_weight[177][38],
reservoir_weight[177][39],
reservoir_weight[177][40],
reservoir_weight[177][41],
reservoir_weight[177][42],
reservoir_weight[177][43],
reservoir_weight[177][44],
reservoir_weight[177][45],
reservoir_weight[177][46],
reservoir_weight[177][47],
reservoir_weight[177][48],
reservoir_weight[177][49],
reservoir_weight[177][50],
reservoir_weight[177][51],
reservoir_weight[177][52],
reservoir_weight[177][53],
reservoir_weight[177][54],
reservoir_weight[177][55],
reservoir_weight[177][56],
reservoir_weight[177][57],
reservoir_weight[177][58],
reservoir_weight[177][59],
reservoir_weight[177][60],
reservoir_weight[177][61],
reservoir_weight[177][62],
reservoir_weight[177][63],
reservoir_weight[177][64],
reservoir_weight[177][65],
reservoir_weight[177][66],
reservoir_weight[177][67],
reservoir_weight[177][68],
reservoir_weight[177][69],
reservoir_weight[177][70],
reservoir_weight[177][71],
reservoir_weight[177][72],
reservoir_weight[177][73],
reservoir_weight[177][74],
reservoir_weight[177][75],
reservoir_weight[177][76],
reservoir_weight[177][77],
reservoir_weight[177][78],
reservoir_weight[177][79],
reservoir_weight[177][80],
reservoir_weight[177][81],
reservoir_weight[177][82],
reservoir_weight[177][83],
reservoir_weight[177][84],
reservoir_weight[177][85],
reservoir_weight[177][86],
reservoir_weight[177][87],
reservoir_weight[177][88],
reservoir_weight[177][89],
reservoir_weight[177][90],
reservoir_weight[177][91],
reservoir_weight[177][92],
reservoir_weight[177][93],
reservoir_weight[177][94],
reservoir_weight[177][95],
reservoir_weight[177][96],
reservoir_weight[177][97],
reservoir_weight[177][98],
reservoir_weight[177][99],
reservoir_weight[177][100],
reservoir_weight[177][101],
reservoir_weight[177][102],
reservoir_weight[177][103],
reservoir_weight[177][104],
reservoir_weight[177][105],
reservoir_weight[177][106],
reservoir_weight[177][107],
reservoir_weight[177][108],
reservoir_weight[177][109],
reservoir_weight[177][110],
reservoir_weight[177][111],
reservoir_weight[177][112],
reservoir_weight[177][113],
reservoir_weight[177][114],
reservoir_weight[177][115],
reservoir_weight[177][116],
reservoir_weight[177][117],
reservoir_weight[177][118],
reservoir_weight[177][119],
reservoir_weight[177][120],
reservoir_weight[177][121],
reservoir_weight[177][122],
reservoir_weight[177][123],
reservoir_weight[177][124],
reservoir_weight[177][125],
reservoir_weight[177][126],
reservoir_weight[177][127],
reservoir_weight[177][128],
reservoir_weight[177][129],
reservoir_weight[177][130],
reservoir_weight[177][131],
reservoir_weight[177][132],
reservoir_weight[177][133],
reservoir_weight[177][134],
reservoir_weight[177][135],
reservoir_weight[177][136],
reservoir_weight[177][137],
reservoir_weight[177][138],
reservoir_weight[177][139],
reservoir_weight[177][140],
reservoir_weight[177][141],
reservoir_weight[177][142],
reservoir_weight[177][143],
reservoir_weight[177][144],
reservoir_weight[177][145],
reservoir_weight[177][146],
reservoir_weight[177][147],
reservoir_weight[177][148],
reservoir_weight[177][149],
reservoir_weight[177][150],
reservoir_weight[177][151],
reservoir_weight[177][152],
reservoir_weight[177][153],
reservoir_weight[177][154],
reservoir_weight[177][155],
reservoir_weight[177][156],
reservoir_weight[177][157],
reservoir_weight[177][158],
reservoir_weight[177][159],
reservoir_weight[177][160],
reservoir_weight[177][161],
reservoir_weight[177][162],
reservoir_weight[177][163],
reservoir_weight[177][164],
reservoir_weight[177][165],
reservoir_weight[177][166],
reservoir_weight[177][167],
reservoir_weight[177][168],
reservoir_weight[177][169],
reservoir_weight[177][170],
reservoir_weight[177][171],
reservoir_weight[177][172],
reservoir_weight[177][173],
reservoir_weight[177][174],
reservoir_weight[177][175],
reservoir_weight[177][176],
reservoir_weight[177][177],
reservoir_weight[177][178],
reservoir_weight[177][179],
reservoir_weight[177][180],
reservoir_weight[177][181],
reservoir_weight[177][182],
reservoir_weight[177][183],
reservoir_weight[177][184],
reservoir_weight[177][185],
reservoir_weight[177][186],
reservoir_weight[177][187],
reservoir_weight[177][188],
reservoir_weight[177][189],
reservoir_weight[177][190],
reservoir_weight[177][191],
reservoir_weight[177][192],
reservoir_weight[177][193],
reservoir_weight[177][194],
reservoir_weight[177][195],
reservoir_weight[177][196],
reservoir_weight[177][197],
reservoir_weight[177][198],
reservoir_weight[177][199]
},
{reservoir_weight[178][0],
reservoir_weight[178][1],
reservoir_weight[178][2],
reservoir_weight[178][3],
reservoir_weight[178][4],
reservoir_weight[178][5],
reservoir_weight[178][6],
reservoir_weight[178][7],
reservoir_weight[178][8],
reservoir_weight[178][9],
reservoir_weight[178][10],
reservoir_weight[178][11],
reservoir_weight[178][12],
reservoir_weight[178][13],
reservoir_weight[178][14],
reservoir_weight[178][15],
reservoir_weight[178][16],
reservoir_weight[178][17],
reservoir_weight[178][18],
reservoir_weight[178][19],
reservoir_weight[178][20],
reservoir_weight[178][21],
reservoir_weight[178][22],
reservoir_weight[178][23],
reservoir_weight[178][24],
reservoir_weight[178][25],
reservoir_weight[178][26],
reservoir_weight[178][27],
reservoir_weight[178][28],
reservoir_weight[178][29],
reservoir_weight[178][30],
reservoir_weight[178][31],
reservoir_weight[178][32],
reservoir_weight[178][33],
reservoir_weight[178][34],
reservoir_weight[178][35],
reservoir_weight[178][36],
reservoir_weight[178][37],
reservoir_weight[178][38],
reservoir_weight[178][39],
reservoir_weight[178][40],
reservoir_weight[178][41],
reservoir_weight[178][42],
reservoir_weight[178][43],
reservoir_weight[178][44],
reservoir_weight[178][45],
reservoir_weight[178][46],
reservoir_weight[178][47],
reservoir_weight[178][48],
reservoir_weight[178][49],
reservoir_weight[178][50],
reservoir_weight[178][51],
reservoir_weight[178][52],
reservoir_weight[178][53],
reservoir_weight[178][54],
reservoir_weight[178][55],
reservoir_weight[178][56],
reservoir_weight[178][57],
reservoir_weight[178][58],
reservoir_weight[178][59],
reservoir_weight[178][60],
reservoir_weight[178][61],
reservoir_weight[178][62],
reservoir_weight[178][63],
reservoir_weight[178][64],
reservoir_weight[178][65],
reservoir_weight[178][66],
reservoir_weight[178][67],
reservoir_weight[178][68],
reservoir_weight[178][69],
reservoir_weight[178][70],
reservoir_weight[178][71],
reservoir_weight[178][72],
reservoir_weight[178][73],
reservoir_weight[178][74],
reservoir_weight[178][75],
reservoir_weight[178][76],
reservoir_weight[178][77],
reservoir_weight[178][78],
reservoir_weight[178][79],
reservoir_weight[178][80],
reservoir_weight[178][81],
reservoir_weight[178][82],
reservoir_weight[178][83],
reservoir_weight[178][84],
reservoir_weight[178][85],
reservoir_weight[178][86],
reservoir_weight[178][87],
reservoir_weight[178][88],
reservoir_weight[178][89],
reservoir_weight[178][90],
reservoir_weight[178][91],
reservoir_weight[178][92],
reservoir_weight[178][93],
reservoir_weight[178][94],
reservoir_weight[178][95],
reservoir_weight[178][96],
reservoir_weight[178][97],
reservoir_weight[178][98],
reservoir_weight[178][99],
reservoir_weight[178][100],
reservoir_weight[178][101],
reservoir_weight[178][102],
reservoir_weight[178][103],
reservoir_weight[178][104],
reservoir_weight[178][105],
reservoir_weight[178][106],
reservoir_weight[178][107],
reservoir_weight[178][108],
reservoir_weight[178][109],
reservoir_weight[178][110],
reservoir_weight[178][111],
reservoir_weight[178][112],
reservoir_weight[178][113],
reservoir_weight[178][114],
reservoir_weight[178][115],
reservoir_weight[178][116],
reservoir_weight[178][117],
reservoir_weight[178][118],
reservoir_weight[178][119],
reservoir_weight[178][120],
reservoir_weight[178][121],
reservoir_weight[178][122],
reservoir_weight[178][123],
reservoir_weight[178][124],
reservoir_weight[178][125],
reservoir_weight[178][126],
reservoir_weight[178][127],
reservoir_weight[178][128],
reservoir_weight[178][129],
reservoir_weight[178][130],
reservoir_weight[178][131],
reservoir_weight[178][132],
reservoir_weight[178][133],
reservoir_weight[178][134],
reservoir_weight[178][135],
reservoir_weight[178][136],
reservoir_weight[178][137],
reservoir_weight[178][138],
reservoir_weight[178][139],
reservoir_weight[178][140],
reservoir_weight[178][141],
reservoir_weight[178][142],
reservoir_weight[178][143],
reservoir_weight[178][144],
reservoir_weight[178][145],
reservoir_weight[178][146],
reservoir_weight[178][147],
reservoir_weight[178][148],
reservoir_weight[178][149],
reservoir_weight[178][150],
reservoir_weight[178][151],
reservoir_weight[178][152],
reservoir_weight[178][153],
reservoir_weight[178][154],
reservoir_weight[178][155],
reservoir_weight[178][156],
reservoir_weight[178][157],
reservoir_weight[178][158],
reservoir_weight[178][159],
reservoir_weight[178][160],
reservoir_weight[178][161],
reservoir_weight[178][162],
reservoir_weight[178][163],
reservoir_weight[178][164],
reservoir_weight[178][165],
reservoir_weight[178][166],
reservoir_weight[178][167],
reservoir_weight[178][168],
reservoir_weight[178][169],
reservoir_weight[178][170],
reservoir_weight[178][171],
reservoir_weight[178][172],
reservoir_weight[178][173],
reservoir_weight[178][174],
reservoir_weight[178][175],
reservoir_weight[178][176],
reservoir_weight[178][177],
reservoir_weight[178][178],
reservoir_weight[178][179],
reservoir_weight[178][180],
reservoir_weight[178][181],
reservoir_weight[178][182],
reservoir_weight[178][183],
reservoir_weight[178][184],
reservoir_weight[178][185],
reservoir_weight[178][186],
reservoir_weight[178][187],
reservoir_weight[178][188],
reservoir_weight[178][189],
reservoir_weight[178][190],
reservoir_weight[178][191],
reservoir_weight[178][192],
reservoir_weight[178][193],
reservoir_weight[178][194],
reservoir_weight[178][195],
reservoir_weight[178][196],
reservoir_weight[178][197],
reservoir_weight[178][198],
reservoir_weight[178][199]
},
{reservoir_weight[179][0],
reservoir_weight[179][1],
reservoir_weight[179][2],
reservoir_weight[179][3],
reservoir_weight[179][4],
reservoir_weight[179][5],
reservoir_weight[179][6],
reservoir_weight[179][7],
reservoir_weight[179][8],
reservoir_weight[179][9],
reservoir_weight[179][10],
reservoir_weight[179][11],
reservoir_weight[179][12],
reservoir_weight[179][13],
reservoir_weight[179][14],
reservoir_weight[179][15],
reservoir_weight[179][16],
reservoir_weight[179][17],
reservoir_weight[179][18],
reservoir_weight[179][19],
reservoir_weight[179][20],
reservoir_weight[179][21],
reservoir_weight[179][22],
reservoir_weight[179][23],
reservoir_weight[179][24],
reservoir_weight[179][25],
reservoir_weight[179][26],
reservoir_weight[179][27],
reservoir_weight[179][28],
reservoir_weight[179][29],
reservoir_weight[179][30],
reservoir_weight[179][31],
reservoir_weight[179][32],
reservoir_weight[179][33],
reservoir_weight[179][34],
reservoir_weight[179][35],
reservoir_weight[179][36],
reservoir_weight[179][37],
reservoir_weight[179][38],
reservoir_weight[179][39],
reservoir_weight[179][40],
reservoir_weight[179][41],
reservoir_weight[179][42],
reservoir_weight[179][43],
reservoir_weight[179][44],
reservoir_weight[179][45],
reservoir_weight[179][46],
reservoir_weight[179][47],
reservoir_weight[179][48],
reservoir_weight[179][49],
reservoir_weight[179][50],
reservoir_weight[179][51],
reservoir_weight[179][52],
reservoir_weight[179][53],
reservoir_weight[179][54],
reservoir_weight[179][55],
reservoir_weight[179][56],
reservoir_weight[179][57],
reservoir_weight[179][58],
reservoir_weight[179][59],
reservoir_weight[179][60],
reservoir_weight[179][61],
reservoir_weight[179][62],
reservoir_weight[179][63],
reservoir_weight[179][64],
reservoir_weight[179][65],
reservoir_weight[179][66],
reservoir_weight[179][67],
reservoir_weight[179][68],
reservoir_weight[179][69],
reservoir_weight[179][70],
reservoir_weight[179][71],
reservoir_weight[179][72],
reservoir_weight[179][73],
reservoir_weight[179][74],
reservoir_weight[179][75],
reservoir_weight[179][76],
reservoir_weight[179][77],
reservoir_weight[179][78],
reservoir_weight[179][79],
reservoir_weight[179][80],
reservoir_weight[179][81],
reservoir_weight[179][82],
reservoir_weight[179][83],
reservoir_weight[179][84],
reservoir_weight[179][85],
reservoir_weight[179][86],
reservoir_weight[179][87],
reservoir_weight[179][88],
reservoir_weight[179][89],
reservoir_weight[179][90],
reservoir_weight[179][91],
reservoir_weight[179][92],
reservoir_weight[179][93],
reservoir_weight[179][94],
reservoir_weight[179][95],
reservoir_weight[179][96],
reservoir_weight[179][97],
reservoir_weight[179][98],
reservoir_weight[179][99],
reservoir_weight[179][100],
reservoir_weight[179][101],
reservoir_weight[179][102],
reservoir_weight[179][103],
reservoir_weight[179][104],
reservoir_weight[179][105],
reservoir_weight[179][106],
reservoir_weight[179][107],
reservoir_weight[179][108],
reservoir_weight[179][109],
reservoir_weight[179][110],
reservoir_weight[179][111],
reservoir_weight[179][112],
reservoir_weight[179][113],
reservoir_weight[179][114],
reservoir_weight[179][115],
reservoir_weight[179][116],
reservoir_weight[179][117],
reservoir_weight[179][118],
reservoir_weight[179][119],
reservoir_weight[179][120],
reservoir_weight[179][121],
reservoir_weight[179][122],
reservoir_weight[179][123],
reservoir_weight[179][124],
reservoir_weight[179][125],
reservoir_weight[179][126],
reservoir_weight[179][127],
reservoir_weight[179][128],
reservoir_weight[179][129],
reservoir_weight[179][130],
reservoir_weight[179][131],
reservoir_weight[179][132],
reservoir_weight[179][133],
reservoir_weight[179][134],
reservoir_weight[179][135],
reservoir_weight[179][136],
reservoir_weight[179][137],
reservoir_weight[179][138],
reservoir_weight[179][139],
reservoir_weight[179][140],
reservoir_weight[179][141],
reservoir_weight[179][142],
reservoir_weight[179][143],
reservoir_weight[179][144],
reservoir_weight[179][145],
reservoir_weight[179][146],
reservoir_weight[179][147],
reservoir_weight[179][148],
reservoir_weight[179][149],
reservoir_weight[179][150],
reservoir_weight[179][151],
reservoir_weight[179][152],
reservoir_weight[179][153],
reservoir_weight[179][154],
reservoir_weight[179][155],
reservoir_weight[179][156],
reservoir_weight[179][157],
reservoir_weight[179][158],
reservoir_weight[179][159],
reservoir_weight[179][160],
reservoir_weight[179][161],
reservoir_weight[179][162],
reservoir_weight[179][163],
reservoir_weight[179][164],
reservoir_weight[179][165],
reservoir_weight[179][166],
reservoir_weight[179][167],
reservoir_weight[179][168],
reservoir_weight[179][169],
reservoir_weight[179][170],
reservoir_weight[179][171],
reservoir_weight[179][172],
reservoir_weight[179][173],
reservoir_weight[179][174],
reservoir_weight[179][175],
reservoir_weight[179][176],
reservoir_weight[179][177],
reservoir_weight[179][178],
reservoir_weight[179][179],
reservoir_weight[179][180],
reservoir_weight[179][181],
reservoir_weight[179][182],
reservoir_weight[179][183],
reservoir_weight[179][184],
reservoir_weight[179][185],
reservoir_weight[179][186],
reservoir_weight[179][187],
reservoir_weight[179][188],
reservoir_weight[179][189],
reservoir_weight[179][190],
reservoir_weight[179][191],
reservoir_weight[179][192],
reservoir_weight[179][193],
reservoir_weight[179][194],
reservoir_weight[179][195],
reservoir_weight[179][196],
reservoir_weight[179][197],
reservoir_weight[179][198],
reservoir_weight[179][199]
},
{reservoir_weight[180][0],
reservoir_weight[180][1],
reservoir_weight[180][2],
reservoir_weight[180][3],
reservoir_weight[180][4],
reservoir_weight[180][5],
reservoir_weight[180][6],
reservoir_weight[180][7],
reservoir_weight[180][8],
reservoir_weight[180][9],
reservoir_weight[180][10],
reservoir_weight[180][11],
reservoir_weight[180][12],
reservoir_weight[180][13],
reservoir_weight[180][14],
reservoir_weight[180][15],
reservoir_weight[180][16],
reservoir_weight[180][17],
reservoir_weight[180][18],
reservoir_weight[180][19],
reservoir_weight[180][20],
reservoir_weight[180][21],
reservoir_weight[180][22],
reservoir_weight[180][23],
reservoir_weight[180][24],
reservoir_weight[180][25],
reservoir_weight[180][26],
reservoir_weight[180][27],
reservoir_weight[180][28],
reservoir_weight[180][29],
reservoir_weight[180][30],
reservoir_weight[180][31],
reservoir_weight[180][32],
reservoir_weight[180][33],
reservoir_weight[180][34],
reservoir_weight[180][35],
reservoir_weight[180][36],
reservoir_weight[180][37],
reservoir_weight[180][38],
reservoir_weight[180][39],
reservoir_weight[180][40],
reservoir_weight[180][41],
reservoir_weight[180][42],
reservoir_weight[180][43],
reservoir_weight[180][44],
reservoir_weight[180][45],
reservoir_weight[180][46],
reservoir_weight[180][47],
reservoir_weight[180][48],
reservoir_weight[180][49],
reservoir_weight[180][50],
reservoir_weight[180][51],
reservoir_weight[180][52],
reservoir_weight[180][53],
reservoir_weight[180][54],
reservoir_weight[180][55],
reservoir_weight[180][56],
reservoir_weight[180][57],
reservoir_weight[180][58],
reservoir_weight[180][59],
reservoir_weight[180][60],
reservoir_weight[180][61],
reservoir_weight[180][62],
reservoir_weight[180][63],
reservoir_weight[180][64],
reservoir_weight[180][65],
reservoir_weight[180][66],
reservoir_weight[180][67],
reservoir_weight[180][68],
reservoir_weight[180][69],
reservoir_weight[180][70],
reservoir_weight[180][71],
reservoir_weight[180][72],
reservoir_weight[180][73],
reservoir_weight[180][74],
reservoir_weight[180][75],
reservoir_weight[180][76],
reservoir_weight[180][77],
reservoir_weight[180][78],
reservoir_weight[180][79],
reservoir_weight[180][80],
reservoir_weight[180][81],
reservoir_weight[180][82],
reservoir_weight[180][83],
reservoir_weight[180][84],
reservoir_weight[180][85],
reservoir_weight[180][86],
reservoir_weight[180][87],
reservoir_weight[180][88],
reservoir_weight[180][89],
reservoir_weight[180][90],
reservoir_weight[180][91],
reservoir_weight[180][92],
reservoir_weight[180][93],
reservoir_weight[180][94],
reservoir_weight[180][95],
reservoir_weight[180][96],
reservoir_weight[180][97],
reservoir_weight[180][98],
reservoir_weight[180][99],
reservoir_weight[180][100],
reservoir_weight[180][101],
reservoir_weight[180][102],
reservoir_weight[180][103],
reservoir_weight[180][104],
reservoir_weight[180][105],
reservoir_weight[180][106],
reservoir_weight[180][107],
reservoir_weight[180][108],
reservoir_weight[180][109],
reservoir_weight[180][110],
reservoir_weight[180][111],
reservoir_weight[180][112],
reservoir_weight[180][113],
reservoir_weight[180][114],
reservoir_weight[180][115],
reservoir_weight[180][116],
reservoir_weight[180][117],
reservoir_weight[180][118],
reservoir_weight[180][119],
reservoir_weight[180][120],
reservoir_weight[180][121],
reservoir_weight[180][122],
reservoir_weight[180][123],
reservoir_weight[180][124],
reservoir_weight[180][125],
reservoir_weight[180][126],
reservoir_weight[180][127],
reservoir_weight[180][128],
reservoir_weight[180][129],
reservoir_weight[180][130],
reservoir_weight[180][131],
reservoir_weight[180][132],
reservoir_weight[180][133],
reservoir_weight[180][134],
reservoir_weight[180][135],
reservoir_weight[180][136],
reservoir_weight[180][137],
reservoir_weight[180][138],
reservoir_weight[180][139],
reservoir_weight[180][140],
reservoir_weight[180][141],
reservoir_weight[180][142],
reservoir_weight[180][143],
reservoir_weight[180][144],
reservoir_weight[180][145],
reservoir_weight[180][146],
reservoir_weight[180][147],
reservoir_weight[180][148],
reservoir_weight[180][149],
reservoir_weight[180][150],
reservoir_weight[180][151],
reservoir_weight[180][152],
reservoir_weight[180][153],
reservoir_weight[180][154],
reservoir_weight[180][155],
reservoir_weight[180][156],
reservoir_weight[180][157],
reservoir_weight[180][158],
reservoir_weight[180][159],
reservoir_weight[180][160],
reservoir_weight[180][161],
reservoir_weight[180][162],
reservoir_weight[180][163],
reservoir_weight[180][164],
reservoir_weight[180][165],
reservoir_weight[180][166],
reservoir_weight[180][167],
reservoir_weight[180][168],
reservoir_weight[180][169],
reservoir_weight[180][170],
reservoir_weight[180][171],
reservoir_weight[180][172],
reservoir_weight[180][173],
reservoir_weight[180][174],
reservoir_weight[180][175],
reservoir_weight[180][176],
reservoir_weight[180][177],
reservoir_weight[180][178],
reservoir_weight[180][179],
reservoir_weight[180][180],
reservoir_weight[180][181],
reservoir_weight[180][182],
reservoir_weight[180][183],
reservoir_weight[180][184],
reservoir_weight[180][185],
reservoir_weight[180][186],
reservoir_weight[180][187],
reservoir_weight[180][188],
reservoir_weight[180][189],
reservoir_weight[180][190],
reservoir_weight[180][191],
reservoir_weight[180][192],
reservoir_weight[180][193],
reservoir_weight[180][194],
reservoir_weight[180][195],
reservoir_weight[180][196],
reservoir_weight[180][197],
reservoir_weight[180][198],
reservoir_weight[180][199]
},
{reservoir_weight[181][0],
reservoir_weight[181][1],
reservoir_weight[181][2],
reservoir_weight[181][3],
reservoir_weight[181][4],
reservoir_weight[181][5],
reservoir_weight[181][6],
reservoir_weight[181][7],
reservoir_weight[181][8],
reservoir_weight[181][9],
reservoir_weight[181][10],
reservoir_weight[181][11],
reservoir_weight[181][12],
reservoir_weight[181][13],
reservoir_weight[181][14],
reservoir_weight[181][15],
reservoir_weight[181][16],
reservoir_weight[181][17],
reservoir_weight[181][18],
reservoir_weight[181][19],
reservoir_weight[181][20],
reservoir_weight[181][21],
reservoir_weight[181][22],
reservoir_weight[181][23],
reservoir_weight[181][24],
reservoir_weight[181][25],
reservoir_weight[181][26],
reservoir_weight[181][27],
reservoir_weight[181][28],
reservoir_weight[181][29],
reservoir_weight[181][30],
reservoir_weight[181][31],
reservoir_weight[181][32],
reservoir_weight[181][33],
reservoir_weight[181][34],
reservoir_weight[181][35],
reservoir_weight[181][36],
reservoir_weight[181][37],
reservoir_weight[181][38],
reservoir_weight[181][39],
reservoir_weight[181][40],
reservoir_weight[181][41],
reservoir_weight[181][42],
reservoir_weight[181][43],
reservoir_weight[181][44],
reservoir_weight[181][45],
reservoir_weight[181][46],
reservoir_weight[181][47],
reservoir_weight[181][48],
reservoir_weight[181][49],
reservoir_weight[181][50],
reservoir_weight[181][51],
reservoir_weight[181][52],
reservoir_weight[181][53],
reservoir_weight[181][54],
reservoir_weight[181][55],
reservoir_weight[181][56],
reservoir_weight[181][57],
reservoir_weight[181][58],
reservoir_weight[181][59],
reservoir_weight[181][60],
reservoir_weight[181][61],
reservoir_weight[181][62],
reservoir_weight[181][63],
reservoir_weight[181][64],
reservoir_weight[181][65],
reservoir_weight[181][66],
reservoir_weight[181][67],
reservoir_weight[181][68],
reservoir_weight[181][69],
reservoir_weight[181][70],
reservoir_weight[181][71],
reservoir_weight[181][72],
reservoir_weight[181][73],
reservoir_weight[181][74],
reservoir_weight[181][75],
reservoir_weight[181][76],
reservoir_weight[181][77],
reservoir_weight[181][78],
reservoir_weight[181][79],
reservoir_weight[181][80],
reservoir_weight[181][81],
reservoir_weight[181][82],
reservoir_weight[181][83],
reservoir_weight[181][84],
reservoir_weight[181][85],
reservoir_weight[181][86],
reservoir_weight[181][87],
reservoir_weight[181][88],
reservoir_weight[181][89],
reservoir_weight[181][90],
reservoir_weight[181][91],
reservoir_weight[181][92],
reservoir_weight[181][93],
reservoir_weight[181][94],
reservoir_weight[181][95],
reservoir_weight[181][96],
reservoir_weight[181][97],
reservoir_weight[181][98],
reservoir_weight[181][99],
reservoir_weight[181][100],
reservoir_weight[181][101],
reservoir_weight[181][102],
reservoir_weight[181][103],
reservoir_weight[181][104],
reservoir_weight[181][105],
reservoir_weight[181][106],
reservoir_weight[181][107],
reservoir_weight[181][108],
reservoir_weight[181][109],
reservoir_weight[181][110],
reservoir_weight[181][111],
reservoir_weight[181][112],
reservoir_weight[181][113],
reservoir_weight[181][114],
reservoir_weight[181][115],
reservoir_weight[181][116],
reservoir_weight[181][117],
reservoir_weight[181][118],
reservoir_weight[181][119],
reservoir_weight[181][120],
reservoir_weight[181][121],
reservoir_weight[181][122],
reservoir_weight[181][123],
reservoir_weight[181][124],
reservoir_weight[181][125],
reservoir_weight[181][126],
reservoir_weight[181][127],
reservoir_weight[181][128],
reservoir_weight[181][129],
reservoir_weight[181][130],
reservoir_weight[181][131],
reservoir_weight[181][132],
reservoir_weight[181][133],
reservoir_weight[181][134],
reservoir_weight[181][135],
reservoir_weight[181][136],
reservoir_weight[181][137],
reservoir_weight[181][138],
reservoir_weight[181][139],
reservoir_weight[181][140],
reservoir_weight[181][141],
reservoir_weight[181][142],
reservoir_weight[181][143],
reservoir_weight[181][144],
reservoir_weight[181][145],
reservoir_weight[181][146],
reservoir_weight[181][147],
reservoir_weight[181][148],
reservoir_weight[181][149],
reservoir_weight[181][150],
reservoir_weight[181][151],
reservoir_weight[181][152],
reservoir_weight[181][153],
reservoir_weight[181][154],
reservoir_weight[181][155],
reservoir_weight[181][156],
reservoir_weight[181][157],
reservoir_weight[181][158],
reservoir_weight[181][159],
reservoir_weight[181][160],
reservoir_weight[181][161],
reservoir_weight[181][162],
reservoir_weight[181][163],
reservoir_weight[181][164],
reservoir_weight[181][165],
reservoir_weight[181][166],
reservoir_weight[181][167],
reservoir_weight[181][168],
reservoir_weight[181][169],
reservoir_weight[181][170],
reservoir_weight[181][171],
reservoir_weight[181][172],
reservoir_weight[181][173],
reservoir_weight[181][174],
reservoir_weight[181][175],
reservoir_weight[181][176],
reservoir_weight[181][177],
reservoir_weight[181][178],
reservoir_weight[181][179],
reservoir_weight[181][180],
reservoir_weight[181][181],
reservoir_weight[181][182],
reservoir_weight[181][183],
reservoir_weight[181][184],
reservoir_weight[181][185],
reservoir_weight[181][186],
reservoir_weight[181][187],
reservoir_weight[181][188],
reservoir_weight[181][189],
reservoir_weight[181][190],
reservoir_weight[181][191],
reservoir_weight[181][192],
reservoir_weight[181][193],
reservoir_weight[181][194],
reservoir_weight[181][195],
reservoir_weight[181][196],
reservoir_weight[181][197],
reservoir_weight[181][198],
reservoir_weight[181][199]
},
{reservoir_weight[182][0],
reservoir_weight[182][1],
reservoir_weight[182][2],
reservoir_weight[182][3],
reservoir_weight[182][4],
reservoir_weight[182][5],
reservoir_weight[182][6],
reservoir_weight[182][7],
reservoir_weight[182][8],
reservoir_weight[182][9],
reservoir_weight[182][10],
reservoir_weight[182][11],
reservoir_weight[182][12],
reservoir_weight[182][13],
reservoir_weight[182][14],
reservoir_weight[182][15],
reservoir_weight[182][16],
reservoir_weight[182][17],
reservoir_weight[182][18],
reservoir_weight[182][19],
reservoir_weight[182][20],
reservoir_weight[182][21],
reservoir_weight[182][22],
reservoir_weight[182][23],
reservoir_weight[182][24],
reservoir_weight[182][25],
reservoir_weight[182][26],
reservoir_weight[182][27],
reservoir_weight[182][28],
reservoir_weight[182][29],
reservoir_weight[182][30],
reservoir_weight[182][31],
reservoir_weight[182][32],
reservoir_weight[182][33],
reservoir_weight[182][34],
reservoir_weight[182][35],
reservoir_weight[182][36],
reservoir_weight[182][37],
reservoir_weight[182][38],
reservoir_weight[182][39],
reservoir_weight[182][40],
reservoir_weight[182][41],
reservoir_weight[182][42],
reservoir_weight[182][43],
reservoir_weight[182][44],
reservoir_weight[182][45],
reservoir_weight[182][46],
reservoir_weight[182][47],
reservoir_weight[182][48],
reservoir_weight[182][49],
reservoir_weight[182][50],
reservoir_weight[182][51],
reservoir_weight[182][52],
reservoir_weight[182][53],
reservoir_weight[182][54],
reservoir_weight[182][55],
reservoir_weight[182][56],
reservoir_weight[182][57],
reservoir_weight[182][58],
reservoir_weight[182][59],
reservoir_weight[182][60],
reservoir_weight[182][61],
reservoir_weight[182][62],
reservoir_weight[182][63],
reservoir_weight[182][64],
reservoir_weight[182][65],
reservoir_weight[182][66],
reservoir_weight[182][67],
reservoir_weight[182][68],
reservoir_weight[182][69],
reservoir_weight[182][70],
reservoir_weight[182][71],
reservoir_weight[182][72],
reservoir_weight[182][73],
reservoir_weight[182][74],
reservoir_weight[182][75],
reservoir_weight[182][76],
reservoir_weight[182][77],
reservoir_weight[182][78],
reservoir_weight[182][79],
reservoir_weight[182][80],
reservoir_weight[182][81],
reservoir_weight[182][82],
reservoir_weight[182][83],
reservoir_weight[182][84],
reservoir_weight[182][85],
reservoir_weight[182][86],
reservoir_weight[182][87],
reservoir_weight[182][88],
reservoir_weight[182][89],
reservoir_weight[182][90],
reservoir_weight[182][91],
reservoir_weight[182][92],
reservoir_weight[182][93],
reservoir_weight[182][94],
reservoir_weight[182][95],
reservoir_weight[182][96],
reservoir_weight[182][97],
reservoir_weight[182][98],
reservoir_weight[182][99],
reservoir_weight[182][100],
reservoir_weight[182][101],
reservoir_weight[182][102],
reservoir_weight[182][103],
reservoir_weight[182][104],
reservoir_weight[182][105],
reservoir_weight[182][106],
reservoir_weight[182][107],
reservoir_weight[182][108],
reservoir_weight[182][109],
reservoir_weight[182][110],
reservoir_weight[182][111],
reservoir_weight[182][112],
reservoir_weight[182][113],
reservoir_weight[182][114],
reservoir_weight[182][115],
reservoir_weight[182][116],
reservoir_weight[182][117],
reservoir_weight[182][118],
reservoir_weight[182][119],
reservoir_weight[182][120],
reservoir_weight[182][121],
reservoir_weight[182][122],
reservoir_weight[182][123],
reservoir_weight[182][124],
reservoir_weight[182][125],
reservoir_weight[182][126],
reservoir_weight[182][127],
reservoir_weight[182][128],
reservoir_weight[182][129],
reservoir_weight[182][130],
reservoir_weight[182][131],
reservoir_weight[182][132],
reservoir_weight[182][133],
reservoir_weight[182][134],
reservoir_weight[182][135],
reservoir_weight[182][136],
reservoir_weight[182][137],
reservoir_weight[182][138],
reservoir_weight[182][139],
reservoir_weight[182][140],
reservoir_weight[182][141],
reservoir_weight[182][142],
reservoir_weight[182][143],
reservoir_weight[182][144],
reservoir_weight[182][145],
reservoir_weight[182][146],
reservoir_weight[182][147],
reservoir_weight[182][148],
reservoir_weight[182][149],
reservoir_weight[182][150],
reservoir_weight[182][151],
reservoir_weight[182][152],
reservoir_weight[182][153],
reservoir_weight[182][154],
reservoir_weight[182][155],
reservoir_weight[182][156],
reservoir_weight[182][157],
reservoir_weight[182][158],
reservoir_weight[182][159],
reservoir_weight[182][160],
reservoir_weight[182][161],
reservoir_weight[182][162],
reservoir_weight[182][163],
reservoir_weight[182][164],
reservoir_weight[182][165],
reservoir_weight[182][166],
reservoir_weight[182][167],
reservoir_weight[182][168],
reservoir_weight[182][169],
reservoir_weight[182][170],
reservoir_weight[182][171],
reservoir_weight[182][172],
reservoir_weight[182][173],
reservoir_weight[182][174],
reservoir_weight[182][175],
reservoir_weight[182][176],
reservoir_weight[182][177],
reservoir_weight[182][178],
reservoir_weight[182][179],
reservoir_weight[182][180],
reservoir_weight[182][181],
reservoir_weight[182][182],
reservoir_weight[182][183],
reservoir_weight[182][184],
reservoir_weight[182][185],
reservoir_weight[182][186],
reservoir_weight[182][187],
reservoir_weight[182][188],
reservoir_weight[182][189],
reservoir_weight[182][190],
reservoir_weight[182][191],
reservoir_weight[182][192],
reservoir_weight[182][193],
reservoir_weight[182][194],
reservoir_weight[182][195],
reservoir_weight[182][196],
reservoir_weight[182][197],
reservoir_weight[182][198],
reservoir_weight[182][199]
},
{reservoir_weight[183][0],
reservoir_weight[183][1],
reservoir_weight[183][2],
reservoir_weight[183][3],
reservoir_weight[183][4],
reservoir_weight[183][5],
reservoir_weight[183][6],
reservoir_weight[183][7],
reservoir_weight[183][8],
reservoir_weight[183][9],
reservoir_weight[183][10],
reservoir_weight[183][11],
reservoir_weight[183][12],
reservoir_weight[183][13],
reservoir_weight[183][14],
reservoir_weight[183][15],
reservoir_weight[183][16],
reservoir_weight[183][17],
reservoir_weight[183][18],
reservoir_weight[183][19],
reservoir_weight[183][20],
reservoir_weight[183][21],
reservoir_weight[183][22],
reservoir_weight[183][23],
reservoir_weight[183][24],
reservoir_weight[183][25],
reservoir_weight[183][26],
reservoir_weight[183][27],
reservoir_weight[183][28],
reservoir_weight[183][29],
reservoir_weight[183][30],
reservoir_weight[183][31],
reservoir_weight[183][32],
reservoir_weight[183][33],
reservoir_weight[183][34],
reservoir_weight[183][35],
reservoir_weight[183][36],
reservoir_weight[183][37],
reservoir_weight[183][38],
reservoir_weight[183][39],
reservoir_weight[183][40],
reservoir_weight[183][41],
reservoir_weight[183][42],
reservoir_weight[183][43],
reservoir_weight[183][44],
reservoir_weight[183][45],
reservoir_weight[183][46],
reservoir_weight[183][47],
reservoir_weight[183][48],
reservoir_weight[183][49],
reservoir_weight[183][50],
reservoir_weight[183][51],
reservoir_weight[183][52],
reservoir_weight[183][53],
reservoir_weight[183][54],
reservoir_weight[183][55],
reservoir_weight[183][56],
reservoir_weight[183][57],
reservoir_weight[183][58],
reservoir_weight[183][59],
reservoir_weight[183][60],
reservoir_weight[183][61],
reservoir_weight[183][62],
reservoir_weight[183][63],
reservoir_weight[183][64],
reservoir_weight[183][65],
reservoir_weight[183][66],
reservoir_weight[183][67],
reservoir_weight[183][68],
reservoir_weight[183][69],
reservoir_weight[183][70],
reservoir_weight[183][71],
reservoir_weight[183][72],
reservoir_weight[183][73],
reservoir_weight[183][74],
reservoir_weight[183][75],
reservoir_weight[183][76],
reservoir_weight[183][77],
reservoir_weight[183][78],
reservoir_weight[183][79],
reservoir_weight[183][80],
reservoir_weight[183][81],
reservoir_weight[183][82],
reservoir_weight[183][83],
reservoir_weight[183][84],
reservoir_weight[183][85],
reservoir_weight[183][86],
reservoir_weight[183][87],
reservoir_weight[183][88],
reservoir_weight[183][89],
reservoir_weight[183][90],
reservoir_weight[183][91],
reservoir_weight[183][92],
reservoir_weight[183][93],
reservoir_weight[183][94],
reservoir_weight[183][95],
reservoir_weight[183][96],
reservoir_weight[183][97],
reservoir_weight[183][98],
reservoir_weight[183][99],
reservoir_weight[183][100],
reservoir_weight[183][101],
reservoir_weight[183][102],
reservoir_weight[183][103],
reservoir_weight[183][104],
reservoir_weight[183][105],
reservoir_weight[183][106],
reservoir_weight[183][107],
reservoir_weight[183][108],
reservoir_weight[183][109],
reservoir_weight[183][110],
reservoir_weight[183][111],
reservoir_weight[183][112],
reservoir_weight[183][113],
reservoir_weight[183][114],
reservoir_weight[183][115],
reservoir_weight[183][116],
reservoir_weight[183][117],
reservoir_weight[183][118],
reservoir_weight[183][119],
reservoir_weight[183][120],
reservoir_weight[183][121],
reservoir_weight[183][122],
reservoir_weight[183][123],
reservoir_weight[183][124],
reservoir_weight[183][125],
reservoir_weight[183][126],
reservoir_weight[183][127],
reservoir_weight[183][128],
reservoir_weight[183][129],
reservoir_weight[183][130],
reservoir_weight[183][131],
reservoir_weight[183][132],
reservoir_weight[183][133],
reservoir_weight[183][134],
reservoir_weight[183][135],
reservoir_weight[183][136],
reservoir_weight[183][137],
reservoir_weight[183][138],
reservoir_weight[183][139],
reservoir_weight[183][140],
reservoir_weight[183][141],
reservoir_weight[183][142],
reservoir_weight[183][143],
reservoir_weight[183][144],
reservoir_weight[183][145],
reservoir_weight[183][146],
reservoir_weight[183][147],
reservoir_weight[183][148],
reservoir_weight[183][149],
reservoir_weight[183][150],
reservoir_weight[183][151],
reservoir_weight[183][152],
reservoir_weight[183][153],
reservoir_weight[183][154],
reservoir_weight[183][155],
reservoir_weight[183][156],
reservoir_weight[183][157],
reservoir_weight[183][158],
reservoir_weight[183][159],
reservoir_weight[183][160],
reservoir_weight[183][161],
reservoir_weight[183][162],
reservoir_weight[183][163],
reservoir_weight[183][164],
reservoir_weight[183][165],
reservoir_weight[183][166],
reservoir_weight[183][167],
reservoir_weight[183][168],
reservoir_weight[183][169],
reservoir_weight[183][170],
reservoir_weight[183][171],
reservoir_weight[183][172],
reservoir_weight[183][173],
reservoir_weight[183][174],
reservoir_weight[183][175],
reservoir_weight[183][176],
reservoir_weight[183][177],
reservoir_weight[183][178],
reservoir_weight[183][179],
reservoir_weight[183][180],
reservoir_weight[183][181],
reservoir_weight[183][182],
reservoir_weight[183][183],
reservoir_weight[183][184],
reservoir_weight[183][185],
reservoir_weight[183][186],
reservoir_weight[183][187],
reservoir_weight[183][188],
reservoir_weight[183][189],
reservoir_weight[183][190],
reservoir_weight[183][191],
reservoir_weight[183][192],
reservoir_weight[183][193],
reservoir_weight[183][194],
reservoir_weight[183][195],
reservoir_weight[183][196],
reservoir_weight[183][197],
reservoir_weight[183][198],
reservoir_weight[183][199]
},
{reservoir_weight[184][0],
reservoir_weight[184][1],
reservoir_weight[184][2],
reservoir_weight[184][3],
reservoir_weight[184][4],
reservoir_weight[184][5],
reservoir_weight[184][6],
reservoir_weight[184][7],
reservoir_weight[184][8],
reservoir_weight[184][9],
reservoir_weight[184][10],
reservoir_weight[184][11],
reservoir_weight[184][12],
reservoir_weight[184][13],
reservoir_weight[184][14],
reservoir_weight[184][15],
reservoir_weight[184][16],
reservoir_weight[184][17],
reservoir_weight[184][18],
reservoir_weight[184][19],
reservoir_weight[184][20],
reservoir_weight[184][21],
reservoir_weight[184][22],
reservoir_weight[184][23],
reservoir_weight[184][24],
reservoir_weight[184][25],
reservoir_weight[184][26],
reservoir_weight[184][27],
reservoir_weight[184][28],
reservoir_weight[184][29],
reservoir_weight[184][30],
reservoir_weight[184][31],
reservoir_weight[184][32],
reservoir_weight[184][33],
reservoir_weight[184][34],
reservoir_weight[184][35],
reservoir_weight[184][36],
reservoir_weight[184][37],
reservoir_weight[184][38],
reservoir_weight[184][39],
reservoir_weight[184][40],
reservoir_weight[184][41],
reservoir_weight[184][42],
reservoir_weight[184][43],
reservoir_weight[184][44],
reservoir_weight[184][45],
reservoir_weight[184][46],
reservoir_weight[184][47],
reservoir_weight[184][48],
reservoir_weight[184][49],
reservoir_weight[184][50],
reservoir_weight[184][51],
reservoir_weight[184][52],
reservoir_weight[184][53],
reservoir_weight[184][54],
reservoir_weight[184][55],
reservoir_weight[184][56],
reservoir_weight[184][57],
reservoir_weight[184][58],
reservoir_weight[184][59],
reservoir_weight[184][60],
reservoir_weight[184][61],
reservoir_weight[184][62],
reservoir_weight[184][63],
reservoir_weight[184][64],
reservoir_weight[184][65],
reservoir_weight[184][66],
reservoir_weight[184][67],
reservoir_weight[184][68],
reservoir_weight[184][69],
reservoir_weight[184][70],
reservoir_weight[184][71],
reservoir_weight[184][72],
reservoir_weight[184][73],
reservoir_weight[184][74],
reservoir_weight[184][75],
reservoir_weight[184][76],
reservoir_weight[184][77],
reservoir_weight[184][78],
reservoir_weight[184][79],
reservoir_weight[184][80],
reservoir_weight[184][81],
reservoir_weight[184][82],
reservoir_weight[184][83],
reservoir_weight[184][84],
reservoir_weight[184][85],
reservoir_weight[184][86],
reservoir_weight[184][87],
reservoir_weight[184][88],
reservoir_weight[184][89],
reservoir_weight[184][90],
reservoir_weight[184][91],
reservoir_weight[184][92],
reservoir_weight[184][93],
reservoir_weight[184][94],
reservoir_weight[184][95],
reservoir_weight[184][96],
reservoir_weight[184][97],
reservoir_weight[184][98],
reservoir_weight[184][99],
reservoir_weight[184][100],
reservoir_weight[184][101],
reservoir_weight[184][102],
reservoir_weight[184][103],
reservoir_weight[184][104],
reservoir_weight[184][105],
reservoir_weight[184][106],
reservoir_weight[184][107],
reservoir_weight[184][108],
reservoir_weight[184][109],
reservoir_weight[184][110],
reservoir_weight[184][111],
reservoir_weight[184][112],
reservoir_weight[184][113],
reservoir_weight[184][114],
reservoir_weight[184][115],
reservoir_weight[184][116],
reservoir_weight[184][117],
reservoir_weight[184][118],
reservoir_weight[184][119],
reservoir_weight[184][120],
reservoir_weight[184][121],
reservoir_weight[184][122],
reservoir_weight[184][123],
reservoir_weight[184][124],
reservoir_weight[184][125],
reservoir_weight[184][126],
reservoir_weight[184][127],
reservoir_weight[184][128],
reservoir_weight[184][129],
reservoir_weight[184][130],
reservoir_weight[184][131],
reservoir_weight[184][132],
reservoir_weight[184][133],
reservoir_weight[184][134],
reservoir_weight[184][135],
reservoir_weight[184][136],
reservoir_weight[184][137],
reservoir_weight[184][138],
reservoir_weight[184][139],
reservoir_weight[184][140],
reservoir_weight[184][141],
reservoir_weight[184][142],
reservoir_weight[184][143],
reservoir_weight[184][144],
reservoir_weight[184][145],
reservoir_weight[184][146],
reservoir_weight[184][147],
reservoir_weight[184][148],
reservoir_weight[184][149],
reservoir_weight[184][150],
reservoir_weight[184][151],
reservoir_weight[184][152],
reservoir_weight[184][153],
reservoir_weight[184][154],
reservoir_weight[184][155],
reservoir_weight[184][156],
reservoir_weight[184][157],
reservoir_weight[184][158],
reservoir_weight[184][159],
reservoir_weight[184][160],
reservoir_weight[184][161],
reservoir_weight[184][162],
reservoir_weight[184][163],
reservoir_weight[184][164],
reservoir_weight[184][165],
reservoir_weight[184][166],
reservoir_weight[184][167],
reservoir_weight[184][168],
reservoir_weight[184][169],
reservoir_weight[184][170],
reservoir_weight[184][171],
reservoir_weight[184][172],
reservoir_weight[184][173],
reservoir_weight[184][174],
reservoir_weight[184][175],
reservoir_weight[184][176],
reservoir_weight[184][177],
reservoir_weight[184][178],
reservoir_weight[184][179],
reservoir_weight[184][180],
reservoir_weight[184][181],
reservoir_weight[184][182],
reservoir_weight[184][183],
reservoir_weight[184][184],
reservoir_weight[184][185],
reservoir_weight[184][186],
reservoir_weight[184][187],
reservoir_weight[184][188],
reservoir_weight[184][189],
reservoir_weight[184][190],
reservoir_weight[184][191],
reservoir_weight[184][192],
reservoir_weight[184][193],
reservoir_weight[184][194],
reservoir_weight[184][195],
reservoir_weight[184][196],
reservoir_weight[184][197],
reservoir_weight[184][198],
reservoir_weight[184][199]
},
{reservoir_weight[185][0],
reservoir_weight[185][1],
reservoir_weight[185][2],
reservoir_weight[185][3],
reservoir_weight[185][4],
reservoir_weight[185][5],
reservoir_weight[185][6],
reservoir_weight[185][7],
reservoir_weight[185][8],
reservoir_weight[185][9],
reservoir_weight[185][10],
reservoir_weight[185][11],
reservoir_weight[185][12],
reservoir_weight[185][13],
reservoir_weight[185][14],
reservoir_weight[185][15],
reservoir_weight[185][16],
reservoir_weight[185][17],
reservoir_weight[185][18],
reservoir_weight[185][19],
reservoir_weight[185][20],
reservoir_weight[185][21],
reservoir_weight[185][22],
reservoir_weight[185][23],
reservoir_weight[185][24],
reservoir_weight[185][25],
reservoir_weight[185][26],
reservoir_weight[185][27],
reservoir_weight[185][28],
reservoir_weight[185][29],
reservoir_weight[185][30],
reservoir_weight[185][31],
reservoir_weight[185][32],
reservoir_weight[185][33],
reservoir_weight[185][34],
reservoir_weight[185][35],
reservoir_weight[185][36],
reservoir_weight[185][37],
reservoir_weight[185][38],
reservoir_weight[185][39],
reservoir_weight[185][40],
reservoir_weight[185][41],
reservoir_weight[185][42],
reservoir_weight[185][43],
reservoir_weight[185][44],
reservoir_weight[185][45],
reservoir_weight[185][46],
reservoir_weight[185][47],
reservoir_weight[185][48],
reservoir_weight[185][49],
reservoir_weight[185][50],
reservoir_weight[185][51],
reservoir_weight[185][52],
reservoir_weight[185][53],
reservoir_weight[185][54],
reservoir_weight[185][55],
reservoir_weight[185][56],
reservoir_weight[185][57],
reservoir_weight[185][58],
reservoir_weight[185][59],
reservoir_weight[185][60],
reservoir_weight[185][61],
reservoir_weight[185][62],
reservoir_weight[185][63],
reservoir_weight[185][64],
reservoir_weight[185][65],
reservoir_weight[185][66],
reservoir_weight[185][67],
reservoir_weight[185][68],
reservoir_weight[185][69],
reservoir_weight[185][70],
reservoir_weight[185][71],
reservoir_weight[185][72],
reservoir_weight[185][73],
reservoir_weight[185][74],
reservoir_weight[185][75],
reservoir_weight[185][76],
reservoir_weight[185][77],
reservoir_weight[185][78],
reservoir_weight[185][79],
reservoir_weight[185][80],
reservoir_weight[185][81],
reservoir_weight[185][82],
reservoir_weight[185][83],
reservoir_weight[185][84],
reservoir_weight[185][85],
reservoir_weight[185][86],
reservoir_weight[185][87],
reservoir_weight[185][88],
reservoir_weight[185][89],
reservoir_weight[185][90],
reservoir_weight[185][91],
reservoir_weight[185][92],
reservoir_weight[185][93],
reservoir_weight[185][94],
reservoir_weight[185][95],
reservoir_weight[185][96],
reservoir_weight[185][97],
reservoir_weight[185][98],
reservoir_weight[185][99],
reservoir_weight[185][100],
reservoir_weight[185][101],
reservoir_weight[185][102],
reservoir_weight[185][103],
reservoir_weight[185][104],
reservoir_weight[185][105],
reservoir_weight[185][106],
reservoir_weight[185][107],
reservoir_weight[185][108],
reservoir_weight[185][109],
reservoir_weight[185][110],
reservoir_weight[185][111],
reservoir_weight[185][112],
reservoir_weight[185][113],
reservoir_weight[185][114],
reservoir_weight[185][115],
reservoir_weight[185][116],
reservoir_weight[185][117],
reservoir_weight[185][118],
reservoir_weight[185][119],
reservoir_weight[185][120],
reservoir_weight[185][121],
reservoir_weight[185][122],
reservoir_weight[185][123],
reservoir_weight[185][124],
reservoir_weight[185][125],
reservoir_weight[185][126],
reservoir_weight[185][127],
reservoir_weight[185][128],
reservoir_weight[185][129],
reservoir_weight[185][130],
reservoir_weight[185][131],
reservoir_weight[185][132],
reservoir_weight[185][133],
reservoir_weight[185][134],
reservoir_weight[185][135],
reservoir_weight[185][136],
reservoir_weight[185][137],
reservoir_weight[185][138],
reservoir_weight[185][139],
reservoir_weight[185][140],
reservoir_weight[185][141],
reservoir_weight[185][142],
reservoir_weight[185][143],
reservoir_weight[185][144],
reservoir_weight[185][145],
reservoir_weight[185][146],
reservoir_weight[185][147],
reservoir_weight[185][148],
reservoir_weight[185][149],
reservoir_weight[185][150],
reservoir_weight[185][151],
reservoir_weight[185][152],
reservoir_weight[185][153],
reservoir_weight[185][154],
reservoir_weight[185][155],
reservoir_weight[185][156],
reservoir_weight[185][157],
reservoir_weight[185][158],
reservoir_weight[185][159],
reservoir_weight[185][160],
reservoir_weight[185][161],
reservoir_weight[185][162],
reservoir_weight[185][163],
reservoir_weight[185][164],
reservoir_weight[185][165],
reservoir_weight[185][166],
reservoir_weight[185][167],
reservoir_weight[185][168],
reservoir_weight[185][169],
reservoir_weight[185][170],
reservoir_weight[185][171],
reservoir_weight[185][172],
reservoir_weight[185][173],
reservoir_weight[185][174],
reservoir_weight[185][175],
reservoir_weight[185][176],
reservoir_weight[185][177],
reservoir_weight[185][178],
reservoir_weight[185][179],
reservoir_weight[185][180],
reservoir_weight[185][181],
reservoir_weight[185][182],
reservoir_weight[185][183],
reservoir_weight[185][184],
reservoir_weight[185][185],
reservoir_weight[185][186],
reservoir_weight[185][187],
reservoir_weight[185][188],
reservoir_weight[185][189],
reservoir_weight[185][190],
reservoir_weight[185][191],
reservoir_weight[185][192],
reservoir_weight[185][193],
reservoir_weight[185][194],
reservoir_weight[185][195],
reservoir_weight[185][196],
reservoir_weight[185][197],
reservoir_weight[185][198],
reservoir_weight[185][199]
},
{reservoir_weight[186][0],
reservoir_weight[186][1],
reservoir_weight[186][2],
reservoir_weight[186][3],
reservoir_weight[186][4],
reservoir_weight[186][5],
reservoir_weight[186][6],
reservoir_weight[186][7],
reservoir_weight[186][8],
reservoir_weight[186][9],
reservoir_weight[186][10],
reservoir_weight[186][11],
reservoir_weight[186][12],
reservoir_weight[186][13],
reservoir_weight[186][14],
reservoir_weight[186][15],
reservoir_weight[186][16],
reservoir_weight[186][17],
reservoir_weight[186][18],
reservoir_weight[186][19],
reservoir_weight[186][20],
reservoir_weight[186][21],
reservoir_weight[186][22],
reservoir_weight[186][23],
reservoir_weight[186][24],
reservoir_weight[186][25],
reservoir_weight[186][26],
reservoir_weight[186][27],
reservoir_weight[186][28],
reservoir_weight[186][29],
reservoir_weight[186][30],
reservoir_weight[186][31],
reservoir_weight[186][32],
reservoir_weight[186][33],
reservoir_weight[186][34],
reservoir_weight[186][35],
reservoir_weight[186][36],
reservoir_weight[186][37],
reservoir_weight[186][38],
reservoir_weight[186][39],
reservoir_weight[186][40],
reservoir_weight[186][41],
reservoir_weight[186][42],
reservoir_weight[186][43],
reservoir_weight[186][44],
reservoir_weight[186][45],
reservoir_weight[186][46],
reservoir_weight[186][47],
reservoir_weight[186][48],
reservoir_weight[186][49],
reservoir_weight[186][50],
reservoir_weight[186][51],
reservoir_weight[186][52],
reservoir_weight[186][53],
reservoir_weight[186][54],
reservoir_weight[186][55],
reservoir_weight[186][56],
reservoir_weight[186][57],
reservoir_weight[186][58],
reservoir_weight[186][59],
reservoir_weight[186][60],
reservoir_weight[186][61],
reservoir_weight[186][62],
reservoir_weight[186][63],
reservoir_weight[186][64],
reservoir_weight[186][65],
reservoir_weight[186][66],
reservoir_weight[186][67],
reservoir_weight[186][68],
reservoir_weight[186][69],
reservoir_weight[186][70],
reservoir_weight[186][71],
reservoir_weight[186][72],
reservoir_weight[186][73],
reservoir_weight[186][74],
reservoir_weight[186][75],
reservoir_weight[186][76],
reservoir_weight[186][77],
reservoir_weight[186][78],
reservoir_weight[186][79],
reservoir_weight[186][80],
reservoir_weight[186][81],
reservoir_weight[186][82],
reservoir_weight[186][83],
reservoir_weight[186][84],
reservoir_weight[186][85],
reservoir_weight[186][86],
reservoir_weight[186][87],
reservoir_weight[186][88],
reservoir_weight[186][89],
reservoir_weight[186][90],
reservoir_weight[186][91],
reservoir_weight[186][92],
reservoir_weight[186][93],
reservoir_weight[186][94],
reservoir_weight[186][95],
reservoir_weight[186][96],
reservoir_weight[186][97],
reservoir_weight[186][98],
reservoir_weight[186][99],
reservoir_weight[186][100],
reservoir_weight[186][101],
reservoir_weight[186][102],
reservoir_weight[186][103],
reservoir_weight[186][104],
reservoir_weight[186][105],
reservoir_weight[186][106],
reservoir_weight[186][107],
reservoir_weight[186][108],
reservoir_weight[186][109],
reservoir_weight[186][110],
reservoir_weight[186][111],
reservoir_weight[186][112],
reservoir_weight[186][113],
reservoir_weight[186][114],
reservoir_weight[186][115],
reservoir_weight[186][116],
reservoir_weight[186][117],
reservoir_weight[186][118],
reservoir_weight[186][119],
reservoir_weight[186][120],
reservoir_weight[186][121],
reservoir_weight[186][122],
reservoir_weight[186][123],
reservoir_weight[186][124],
reservoir_weight[186][125],
reservoir_weight[186][126],
reservoir_weight[186][127],
reservoir_weight[186][128],
reservoir_weight[186][129],
reservoir_weight[186][130],
reservoir_weight[186][131],
reservoir_weight[186][132],
reservoir_weight[186][133],
reservoir_weight[186][134],
reservoir_weight[186][135],
reservoir_weight[186][136],
reservoir_weight[186][137],
reservoir_weight[186][138],
reservoir_weight[186][139],
reservoir_weight[186][140],
reservoir_weight[186][141],
reservoir_weight[186][142],
reservoir_weight[186][143],
reservoir_weight[186][144],
reservoir_weight[186][145],
reservoir_weight[186][146],
reservoir_weight[186][147],
reservoir_weight[186][148],
reservoir_weight[186][149],
reservoir_weight[186][150],
reservoir_weight[186][151],
reservoir_weight[186][152],
reservoir_weight[186][153],
reservoir_weight[186][154],
reservoir_weight[186][155],
reservoir_weight[186][156],
reservoir_weight[186][157],
reservoir_weight[186][158],
reservoir_weight[186][159],
reservoir_weight[186][160],
reservoir_weight[186][161],
reservoir_weight[186][162],
reservoir_weight[186][163],
reservoir_weight[186][164],
reservoir_weight[186][165],
reservoir_weight[186][166],
reservoir_weight[186][167],
reservoir_weight[186][168],
reservoir_weight[186][169],
reservoir_weight[186][170],
reservoir_weight[186][171],
reservoir_weight[186][172],
reservoir_weight[186][173],
reservoir_weight[186][174],
reservoir_weight[186][175],
reservoir_weight[186][176],
reservoir_weight[186][177],
reservoir_weight[186][178],
reservoir_weight[186][179],
reservoir_weight[186][180],
reservoir_weight[186][181],
reservoir_weight[186][182],
reservoir_weight[186][183],
reservoir_weight[186][184],
reservoir_weight[186][185],
reservoir_weight[186][186],
reservoir_weight[186][187],
reservoir_weight[186][188],
reservoir_weight[186][189],
reservoir_weight[186][190],
reservoir_weight[186][191],
reservoir_weight[186][192],
reservoir_weight[186][193],
reservoir_weight[186][194],
reservoir_weight[186][195],
reservoir_weight[186][196],
reservoir_weight[186][197],
reservoir_weight[186][198],
reservoir_weight[186][199]
},
{reservoir_weight[187][0],
reservoir_weight[187][1],
reservoir_weight[187][2],
reservoir_weight[187][3],
reservoir_weight[187][4],
reservoir_weight[187][5],
reservoir_weight[187][6],
reservoir_weight[187][7],
reservoir_weight[187][8],
reservoir_weight[187][9],
reservoir_weight[187][10],
reservoir_weight[187][11],
reservoir_weight[187][12],
reservoir_weight[187][13],
reservoir_weight[187][14],
reservoir_weight[187][15],
reservoir_weight[187][16],
reservoir_weight[187][17],
reservoir_weight[187][18],
reservoir_weight[187][19],
reservoir_weight[187][20],
reservoir_weight[187][21],
reservoir_weight[187][22],
reservoir_weight[187][23],
reservoir_weight[187][24],
reservoir_weight[187][25],
reservoir_weight[187][26],
reservoir_weight[187][27],
reservoir_weight[187][28],
reservoir_weight[187][29],
reservoir_weight[187][30],
reservoir_weight[187][31],
reservoir_weight[187][32],
reservoir_weight[187][33],
reservoir_weight[187][34],
reservoir_weight[187][35],
reservoir_weight[187][36],
reservoir_weight[187][37],
reservoir_weight[187][38],
reservoir_weight[187][39],
reservoir_weight[187][40],
reservoir_weight[187][41],
reservoir_weight[187][42],
reservoir_weight[187][43],
reservoir_weight[187][44],
reservoir_weight[187][45],
reservoir_weight[187][46],
reservoir_weight[187][47],
reservoir_weight[187][48],
reservoir_weight[187][49],
reservoir_weight[187][50],
reservoir_weight[187][51],
reservoir_weight[187][52],
reservoir_weight[187][53],
reservoir_weight[187][54],
reservoir_weight[187][55],
reservoir_weight[187][56],
reservoir_weight[187][57],
reservoir_weight[187][58],
reservoir_weight[187][59],
reservoir_weight[187][60],
reservoir_weight[187][61],
reservoir_weight[187][62],
reservoir_weight[187][63],
reservoir_weight[187][64],
reservoir_weight[187][65],
reservoir_weight[187][66],
reservoir_weight[187][67],
reservoir_weight[187][68],
reservoir_weight[187][69],
reservoir_weight[187][70],
reservoir_weight[187][71],
reservoir_weight[187][72],
reservoir_weight[187][73],
reservoir_weight[187][74],
reservoir_weight[187][75],
reservoir_weight[187][76],
reservoir_weight[187][77],
reservoir_weight[187][78],
reservoir_weight[187][79],
reservoir_weight[187][80],
reservoir_weight[187][81],
reservoir_weight[187][82],
reservoir_weight[187][83],
reservoir_weight[187][84],
reservoir_weight[187][85],
reservoir_weight[187][86],
reservoir_weight[187][87],
reservoir_weight[187][88],
reservoir_weight[187][89],
reservoir_weight[187][90],
reservoir_weight[187][91],
reservoir_weight[187][92],
reservoir_weight[187][93],
reservoir_weight[187][94],
reservoir_weight[187][95],
reservoir_weight[187][96],
reservoir_weight[187][97],
reservoir_weight[187][98],
reservoir_weight[187][99],
reservoir_weight[187][100],
reservoir_weight[187][101],
reservoir_weight[187][102],
reservoir_weight[187][103],
reservoir_weight[187][104],
reservoir_weight[187][105],
reservoir_weight[187][106],
reservoir_weight[187][107],
reservoir_weight[187][108],
reservoir_weight[187][109],
reservoir_weight[187][110],
reservoir_weight[187][111],
reservoir_weight[187][112],
reservoir_weight[187][113],
reservoir_weight[187][114],
reservoir_weight[187][115],
reservoir_weight[187][116],
reservoir_weight[187][117],
reservoir_weight[187][118],
reservoir_weight[187][119],
reservoir_weight[187][120],
reservoir_weight[187][121],
reservoir_weight[187][122],
reservoir_weight[187][123],
reservoir_weight[187][124],
reservoir_weight[187][125],
reservoir_weight[187][126],
reservoir_weight[187][127],
reservoir_weight[187][128],
reservoir_weight[187][129],
reservoir_weight[187][130],
reservoir_weight[187][131],
reservoir_weight[187][132],
reservoir_weight[187][133],
reservoir_weight[187][134],
reservoir_weight[187][135],
reservoir_weight[187][136],
reservoir_weight[187][137],
reservoir_weight[187][138],
reservoir_weight[187][139],
reservoir_weight[187][140],
reservoir_weight[187][141],
reservoir_weight[187][142],
reservoir_weight[187][143],
reservoir_weight[187][144],
reservoir_weight[187][145],
reservoir_weight[187][146],
reservoir_weight[187][147],
reservoir_weight[187][148],
reservoir_weight[187][149],
reservoir_weight[187][150],
reservoir_weight[187][151],
reservoir_weight[187][152],
reservoir_weight[187][153],
reservoir_weight[187][154],
reservoir_weight[187][155],
reservoir_weight[187][156],
reservoir_weight[187][157],
reservoir_weight[187][158],
reservoir_weight[187][159],
reservoir_weight[187][160],
reservoir_weight[187][161],
reservoir_weight[187][162],
reservoir_weight[187][163],
reservoir_weight[187][164],
reservoir_weight[187][165],
reservoir_weight[187][166],
reservoir_weight[187][167],
reservoir_weight[187][168],
reservoir_weight[187][169],
reservoir_weight[187][170],
reservoir_weight[187][171],
reservoir_weight[187][172],
reservoir_weight[187][173],
reservoir_weight[187][174],
reservoir_weight[187][175],
reservoir_weight[187][176],
reservoir_weight[187][177],
reservoir_weight[187][178],
reservoir_weight[187][179],
reservoir_weight[187][180],
reservoir_weight[187][181],
reservoir_weight[187][182],
reservoir_weight[187][183],
reservoir_weight[187][184],
reservoir_weight[187][185],
reservoir_weight[187][186],
reservoir_weight[187][187],
reservoir_weight[187][188],
reservoir_weight[187][189],
reservoir_weight[187][190],
reservoir_weight[187][191],
reservoir_weight[187][192],
reservoir_weight[187][193],
reservoir_weight[187][194],
reservoir_weight[187][195],
reservoir_weight[187][196],
reservoir_weight[187][197],
reservoir_weight[187][198],
reservoir_weight[187][199]
},
{reservoir_weight[188][0],
reservoir_weight[188][1],
reservoir_weight[188][2],
reservoir_weight[188][3],
reservoir_weight[188][4],
reservoir_weight[188][5],
reservoir_weight[188][6],
reservoir_weight[188][7],
reservoir_weight[188][8],
reservoir_weight[188][9],
reservoir_weight[188][10],
reservoir_weight[188][11],
reservoir_weight[188][12],
reservoir_weight[188][13],
reservoir_weight[188][14],
reservoir_weight[188][15],
reservoir_weight[188][16],
reservoir_weight[188][17],
reservoir_weight[188][18],
reservoir_weight[188][19],
reservoir_weight[188][20],
reservoir_weight[188][21],
reservoir_weight[188][22],
reservoir_weight[188][23],
reservoir_weight[188][24],
reservoir_weight[188][25],
reservoir_weight[188][26],
reservoir_weight[188][27],
reservoir_weight[188][28],
reservoir_weight[188][29],
reservoir_weight[188][30],
reservoir_weight[188][31],
reservoir_weight[188][32],
reservoir_weight[188][33],
reservoir_weight[188][34],
reservoir_weight[188][35],
reservoir_weight[188][36],
reservoir_weight[188][37],
reservoir_weight[188][38],
reservoir_weight[188][39],
reservoir_weight[188][40],
reservoir_weight[188][41],
reservoir_weight[188][42],
reservoir_weight[188][43],
reservoir_weight[188][44],
reservoir_weight[188][45],
reservoir_weight[188][46],
reservoir_weight[188][47],
reservoir_weight[188][48],
reservoir_weight[188][49],
reservoir_weight[188][50],
reservoir_weight[188][51],
reservoir_weight[188][52],
reservoir_weight[188][53],
reservoir_weight[188][54],
reservoir_weight[188][55],
reservoir_weight[188][56],
reservoir_weight[188][57],
reservoir_weight[188][58],
reservoir_weight[188][59],
reservoir_weight[188][60],
reservoir_weight[188][61],
reservoir_weight[188][62],
reservoir_weight[188][63],
reservoir_weight[188][64],
reservoir_weight[188][65],
reservoir_weight[188][66],
reservoir_weight[188][67],
reservoir_weight[188][68],
reservoir_weight[188][69],
reservoir_weight[188][70],
reservoir_weight[188][71],
reservoir_weight[188][72],
reservoir_weight[188][73],
reservoir_weight[188][74],
reservoir_weight[188][75],
reservoir_weight[188][76],
reservoir_weight[188][77],
reservoir_weight[188][78],
reservoir_weight[188][79],
reservoir_weight[188][80],
reservoir_weight[188][81],
reservoir_weight[188][82],
reservoir_weight[188][83],
reservoir_weight[188][84],
reservoir_weight[188][85],
reservoir_weight[188][86],
reservoir_weight[188][87],
reservoir_weight[188][88],
reservoir_weight[188][89],
reservoir_weight[188][90],
reservoir_weight[188][91],
reservoir_weight[188][92],
reservoir_weight[188][93],
reservoir_weight[188][94],
reservoir_weight[188][95],
reservoir_weight[188][96],
reservoir_weight[188][97],
reservoir_weight[188][98],
reservoir_weight[188][99],
reservoir_weight[188][100],
reservoir_weight[188][101],
reservoir_weight[188][102],
reservoir_weight[188][103],
reservoir_weight[188][104],
reservoir_weight[188][105],
reservoir_weight[188][106],
reservoir_weight[188][107],
reservoir_weight[188][108],
reservoir_weight[188][109],
reservoir_weight[188][110],
reservoir_weight[188][111],
reservoir_weight[188][112],
reservoir_weight[188][113],
reservoir_weight[188][114],
reservoir_weight[188][115],
reservoir_weight[188][116],
reservoir_weight[188][117],
reservoir_weight[188][118],
reservoir_weight[188][119],
reservoir_weight[188][120],
reservoir_weight[188][121],
reservoir_weight[188][122],
reservoir_weight[188][123],
reservoir_weight[188][124],
reservoir_weight[188][125],
reservoir_weight[188][126],
reservoir_weight[188][127],
reservoir_weight[188][128],
reservoir_weight[188][129],
reservoir_weight[188][130],
reservoir_weight[188][131],
reservoir_weight[188][132],
reservoir_weight[188][133],
reservoir_weight[188][134],
reservoir_weight[188][135],
reservoir_weight[188][136],
reservoir_weight[188][137],
reservoir_weight[188][138],
reservoir_weight[188][139],
reservoir_weight[188][140],
reservoir_weight[188][141],
reservoir_weight[188][142],
reservoir_weight[188][143],
reservoir_weight[188][144],
reservoir_weight[188][145],
reservoir_weight[188][146],
reservoir_weight[188][147],
reservoir_weight[188][148],
reservoir_weight[188][149],
reservoir_weight[188][150],
reservoir_weight[188][151],
reservoir_weight[188][152],
reservoir_weight[188][153],
reservoir_weight[188][154],
reservoir_weight[188][155],
reservoir_weight[188][156],
reservoir_weight[188][157],
reservoir_weight[188][158],
reservoir_weight[188][159],
reservoir_weight[188][160],
reservoir_weight[188][161],
reservoir_weight[188][162],
reservoir_weight[188][163],
reservoir_weight[188][164],
reservoir_weight[188][165],
reservoir_weight[188][166],
reservoir_weight[188][167],
reservoir_weight[188][168],
reservoir_weight[188][169],
reservoir_weight[188][170],
reservoir_weight[188][171],
reservoir_weight[188][172],
reservoir_weight[188][173],
reservoir_weight[188][174],
reservoir_weight[188][175],
reservoir_weight[188][176],
reservoir_weight[188][177],
reservoir_weight[188][178],
reservoir_weight[188][179],
reservoir_weight[188][180],
reservoir_weight[188][181],
reservoir_weight[188][182],
reservoir_weight[188][183],
reservoir_weight[188][184],
reservoir_weight[188][185],
reservoir_weight[188][186],
reservoir_weight[188][187],
reservoir_weight[188][188],
reservoir_weight[188][189],
reservoir_weight[188][190],
reservoir_weight[188][191],
reservoir_weight[188][192],
reservoir_weight[188][193],
reservoir_weight[188][194],
reservoir_weight[188][195],
reservoir_weight[188][196],
reservoir_weight[188][197],
reservoir_weight[188][198],
reservoir_weight[188][199]
},
{reservoir_weight[189][0],
reservoir_weight[189][1],
reservoir_weight[189][2],
reservoir_weight[189][3],
reservoir_weight[189][4],
reservoir_weight[189][5],
reservoir_weight[189][6],
reservoir_weight[189][7],
reservoir_weight[189][8],
reservoir_weight[189][9],
reservoir_weight[189][10],
reservoir_weight[189][11],
reservoir_weight[189][12],
reservoir_weight[189][13],
reservoir_weight[189][14],
reservoir_weight[189][15],
reservoir_weight[189][16],
reservoir_weight[189][17],
reservoir_weight[189][18],
reservoir_weight[189][19],
reservoir_weight[189][20],
reservoir_weight[189][21],
reservoir_weight[189][22],
reservoir_weight[189][23],
reservoir_weight[189][24],
reservoir_weight[189][25],
reservoir_weight[189][26],
reservoir_weight[189][27],
reservoir_weight[189][28],
reservoir_weight[189][29],
reservoir_weight[189][30],
reservoir_weight[189][31],
reservoir_weight[189][32],
reservoir_weight[189][33],
reservoir_weight[189][34],
reservoir_weight[189][35],
reservoir_weight[189][36],
reservoir_weight[189][37],
reservoir_weight[189][38],
reservoir_weight[189][39],
reservoir_weight[189][40],
reservoir_weight[189][41],
reservoir_weight[189][42],
reservoir_weight[189][43],
reservoir_weight[189][44],
reservoir_weight[189][45],
reservoir_weight[189][46],
reservoir_weight[189][47],
reservoir_weight[189][48],
reservoir_weight[189][49],
reservoir_weight[189][50],
reservoir_weight[189][51],
reservoir_weight[189][52],
reservoir_weight[189][53],
reservoir_weight[189][54],
reservoir_weight[189][55],
reservoir_weight[189][56],
reservoir_weight[189][57],
reservoir_weight[189][58],
reservoir_weight[189][59],
reservoir_weight[189][60],
reservoir_weight[189][61],
reservoir_weight[189][62],
reservoir_weight[189][63],
reservoir_weight[189][64],
reservoir_weight[189][65],
reservoir_weight[189][66],
reservoir_weight[189][67],
reservoir_weight[189][68],
reservoir_weight[189][69],
reservoir_weight[189][70],
reservoir_weight[189][71],
reservoir_weight[189][72],
reservoir_weight[189][73],
reservoir_weight[189][74],
reservoir_weight[189][75],
reservoir_weight[189][76],
reservoir_weight[189][77],
reservoir_weight[189][78],
reservoir_weight[189][79],
reservoir_weight[189][80],
reservoir_weight[189][81],
reservoir_weight[189][82],
reservoir_weight[189][83],
reservoir_weight[189][84],
reservoir_weight[189][85],
reservoir_weight[189][86],
reservoir_weight[189][87],
reservoir_weight[189][88],
reservoir_weight[189][89],
reservoir_weight[189][90],
reservoir_weight[189][91],
reservoir_weight[189][92],
reservoir_weight[189][93],
reservoir_weight[189][94],
reservoir_weight[189][95],
reservoir_weight[189][96],
reservoir_weight[189][97],
reservoir_weight[189][98],
reservoir_weight[189][99],
reservoir_weight[189][100],
reservoir_weight[189][101],
reservoir_weight[189][102],
reservoir_weight[189][103],
reservoir_weight[189][104],
reservoir_weight[189][105],
reservoir_weight[189][106],
reservoir_weight[189][107],
reservoir_weight[189][108],
reservoir_weight[189][109],
reservoir_weight[189][110],
reservoir_weight[189][111],
reservoir_weight[189][112],
reservoir_weight[189][113],
reservoir_weight[189][114],
reservoir_weight[189][115],
reservoir_weight[189][116],
reservoir_weight[189][117],
reservoir_weight[189][118],
reservoir_weight[189][119],
reservoir_weight[189][120],
reservoir_weight[189][121],
reservoir_weight[189][122],
reservoir_weight[189][123],
reservoir_weight[189][124],
reservoir_weight[189][125],
reservoir_weight[189][126],
reservoir_weight[189][127],
reservoir_weight[189][128],
reservoir_weight[189][129],
reservoir_weight[189][130],
reservoir_weight[189][131],
reservoir_weight[189][132],
reservoir_weight[189][133],
reservoir_weight[189][134],
reservoir_weight[189][135],
reservoir_weight[189][136],
reservoir_weight[189][137],
reservoir_weight[189][138],
reservoir_weight[189][139],
reservoir_weight[189][140],
reservoir_weight[189][141],
reservoir_weight[189][142],
reservoir_weight[189][143],
reservoir_weight[189][144],
reservoir_weight[189][145],
reservoir_weight[189][146],
reservoir_weight[189][147],
reservoir_weight[189][148],
reservoir_weight[189][149],
reservoir_weight[189][150],
reservoir_weight[189][151],
reservoir_weight[189][152],
reservoir_weight[189][153],
reservoir_weight[189][154],
reservoir_weight[189][155],
reservoir_weight[189][156],
reservoir_weight[189][157],
reservoir_weight[189][158],
reservoir_weight[189][159],
reservoir_weight[189][160],
reservoir_weight[189][161],
reservoir_weight[189][162],
reservoir_weight[189][163],
reservoir_weight[189][164],
reservoir_weight[189][165],
reservoir_weight[189][166],
reservoir_weight[189][167],
reservoir_weight[189][168],
reservoir_weight[189][169],
reservoir_weight[189][170],
reservoir_weight[189][171],
reservoir_weight[189][172],
reservoir_weight[189][173],
reservoir_weight[189][174],
reservoir_weight[189][175],
reservoir_weight[189][176],
reservoir_weight[189][177],
reservoir_weight[189][178],
reservoir_weight[189][179],
reservoir_weight[189][180],
reservoir_weight[189][181],
reservoir_weight[189][182],
reservoir_weight[189][183],
reservoir_weight[189][184],
reservoir_weight[189][185],
reservoir_weight[189][186],
reservoir_weight[189][187],
reservoir_weight[189][188],
reservoir_weight[189][189],
reservoir_weight[189][190],
reservoir_weight[189][191],
reservoir_weight[189][192],
reservoir_weight[189][193],
reservoir_weight[189][194],
reservoir_weight[189][195],
reservoir_weight[189][196],
reservoir_weight[189][197],
reservoir_weight[189][198],
reservoir_weight[189][199]
},
{reservoir_weight[190][0],
reservoir_weight[190][1],
reservoir_weight[190][2],
reservoir_weight[190][3],
reservoir_weight[190][4],
reservoir_weight[190][5],
reservoir_weight[190][6],
reservoir_weight[190][7],
reservoir_weight[190][8],
reservoir_weight[190][9],
reservoir_weight[190][10],
reservoir_weight[190][11],
reservoir_weight[190][12],
reservoir_weight[190][13],
reservoir_weight[190][14],
reservoir_weight[190][15],
reservoir_weight[190][16],
reservoir_weight[190][17],
reservoir_weight[190][18],
reservoir_weight[190][19],
reservoir_weight[190][20],
reservoir_weight[190][21],
reservoir_weight[190][22],
reservoir_weight[190][23],
reservoir_weight[190][24],
reservoir_weight[190][25],
reservoir_weight[190][26],
reservoir_weight[190][27],
reservoir_weight[190][28],
reservoir_weight[190][29],
reservoir_weight[190][30],
reservoir_weight[190][31],
reservoir_weight[190][32],
reservoir_weight[190][33],
reservoir_weight[190][34],
reservoir_weight[190][35],
reservoir_weight[190][36],
reservoir_weight[190][37],
reservoir_weight[190][38],
reservoir_weight[190][39],
reservoir_weight[190][40],
reservoir_weight[190][41],
reservoir_weight[190][42],
reservoir_weight[190][43],
reservoir_weight[190][44],
reservoir_weight[190][45],
reservoir_weight[190][46],
reservoir_weight[190][47],
reservoir_weight[190][48],
reservoir_weight[190][49],
reservoir_weight[190][50],
reservoir_weight[190][51],
reservoir_weight[190][52],
reservoir_weight[190][53],
reservoir_weight[190][54],
reservoir_weight[190][55],
reservoir_weight[190][56],
reservoir_weight[190][57],
reservoir_weight[190][58],
reservoir_weight[190][59],
reservoir_weight[190][60],
reservoir_weight[190][61],
reservoir_weight[190][62],
reservoir_weight[190][63],
reservoir_weight[190][64],
reservoir_weight[190][65],
reservoir_weight[190][66],
reservoir_weight[190][67],
reservoir_weight[190][68],
reservoir_weight[190][69],
reservoir_weight[190][70],
reservoir_weight[190][71],
reservoir_weight[190][72],
reservoir_weight[190][73],
reservoir_weight[190][74],
reservoir_weight[190][75],
reservoir_weight[190][76],
reservoir_weight[190][77],
reservoir_weight[190][78],
reservoir_weight[190][79],
reservoir_weight[190][80],
reservoir_weight[190][81],
reservoir_weight[190][82],
reservoir_weight[190][83],
reservoir_weight[190][84],
reservoir_weight[190][85],
reservoir_weight[190][86],
reservoir_weight[190][87],
reservoir_weight[190][88],
reservoir_weight[190][89],
reservoir_weight[190][90],
reservoir_weight[190][91],
reservoir_weight[190][92],
reservoir_weight[190][93],
reservoir_weight[190][94],
reservoir_weight[190][95],
reservoir_weight[190][96],
reservoir_weight[190][97],
reservoir_weight[190][98],
reservoir_weight[190][99],
reservoir_weight[190][100],
reservoir_weight[190][101],
reservoir_weight[190][102],
reservoir_weight[190][103],
reservoir_weight[190][104],
reservoir_weight[190][105],
reservoir_weight[190][106],
reservoir_weight[190][107],
reservoir_weight[190][108],
reservoir_weight[190][109],
reservoir_weight[190][110],
reservoir_weight[190][111],
reservoir_weight[190][112],
reservoir_weight[190][113],
reservoir_weight[190][114],
reservoir_weight[190][115],
reservoir_weight[190][116],
reservoir_weight[190][117],
reservoir_weight[190][118],
reservoir_weight[190][119],
reservoir_weight[190][120],
reservoir_weight[190][121],
reservoir_weight[190][122],
reservoir_weight[190][123],
reservoir_weight[190][124],
reservoir_weight[190][125],
reservoir_weight[190][126],
reservoir_weight[190][127],
reservoir_weight[190][128],
reservoir_weight[190][129],
reservoir_weight[190][130],
reservoir_weight[190][131],
reservoir_weight[190][132],
reservoir_weight[190][133],
reservoir_weight[190][134],
reservoir_weight[190][135],
reservoir_weight[190][136],
reservoir_weight[190][137],
reservoir_weight[190][138],
reservoir_weight[190][139],
reservoir_weight[190][140],
reservoir_weight[190][141],
reservoir_weight[190][142],
reservoir_weight[190][143],
reservoir_weight[190][144],
reservoir_weight[190][145],
reservoir_weight[190][146],
reservoir_weight[190][147],
reservoir_weight[190][148],
reservoir_weight[190][149],
reservoir_weight[190][150],
reservoir_weight[190][151],
reservoir_weight[190][152],
reservoir_weight[190][153],
reservoir_weight[190][154],
reservoir_weight[190][155],
reservoir_weight[190][156],
reservoir_weight[190][157],
reservoir_weight[190][158],
reservoir_weight[190][159],
reservoir_weight[190][160],
reservoir_weight[190][161],
reservoir_weight[190][162],
reservoir_weight[190][163],
reservoir_weight[190][164],
reservoir_weight[190][165],
reservoir_weight[190][166],
reservoir_weight[190][167],
reservoir_weight[190][168],
reservoir_weight[190][169],
reservoir_weight[190][170],
reservoir_weight[190][171],
reservoir_weight[190][172],
reservoir_weight[190][173],
reservoir_weight[190][174],
reservoir_weight[190][175],
reservoir_weight[190][176],
reservoir_weight[190][177],
reservoir_weight[190][178],
reservoir_weight[190][179],
reservoir_weight[190][180],
reservoir_weight[190][181],
reservoir_weight[190][182],
reservoir_weight[190][183],
reservoir_weight[190][184],
reservoir_weight[190][185],
reservoir_weight[190][186],
reservoir_weight[190][187],
reservoir_weight[190][188],
reservoir_weight[190][189],
reservoir_weight[190][190],
reservoir_weight[190][191],
reservoir_weight[190][192],
reservoir_weight[190][193],
reservoir_weight[190][194],
reservoir_weight[190][195],
reservoir_weight[190][196],
reservoir_weight[190][197],
reservoir_weight[190][198],
reservoir_weight[190][199]
},
{reservoir_weight[191][0],
reservoir_weight[191][1],
reservoir_weight[191][2],
reservoir_weight[191][3],
reservoir_weight[191][4],
reservoir_weight[191][5],
reservoir_weight[191][6],
reservoir_weight[191][7],
reservoir_weight[191][8],
reservoir_weight[191][9],
reservoir_weight[191][10],
reservoir_weight[191][11],
reservoir_weight[191][12],
reservoir_weight[191][13],
reservoir_weight[191][14],
reservoir_weight[191][15],
reservoir_weight[191][16],
reservoir_weight[191][17],
reservoir_weight[191][18],
reservoir_weight[191][19],
reservoir_weight[191][20],
reservoir_weight[191][21],
reservoir_weight[191][22],
reservoir_weight[191][23],
reservoir_weight[191][24],
reservoir_weight[191][25],
reservoir_weight[191][26],
reservoir_weight[191][27],
reservoir_weight[191][28],
reservoir_weight[191][29],
reservoir_weight[191][30],
reservoir_weight[191][31],
reservoir_weight[191][32],
reservoir_weight[191][33],
reservoir_weight[191][34],
reservoir_weight[191][35],
reservoir_weight[191][36],
reservoir_weight[191][37],
reservoir_weight[191][38],
reservoir_weight[191][39],
reservoir_weight[191][40],
reservoir_weight[191][41],
reservoir_weight[191][42],
reservoir_weight[191][43],
reservoir_weight[191][44],
reservoir_weight[191][45],
reservoir_weight[191][46],
reservoir_weight[191][47],
reservoir_weight[191][48],
reservoir_weight[191][49],
reservoir_weight[191][50],
reservoir_weight[191][51],
reservoir_weight[191][52],
reservoir_weight[191][53],
reservoir_weight[191][54],
reservoir_weight[191][55],
reservoir_weight[191][56],
reservoir_weight[191][57],
reservoir_weight[191][58],
reservoir_weight[191][59],
reservoir_weight[191][60],
reservoir_weight[191][61],
reservoir_weight[191][62],
reservoir_weight[191][63],
reservoir_weight[191][64],
reservoir_weight[191][65],
reservoir_weight[191][66],
reservoir_weight[191][67],
reservoir_weight[191][68],
reservoir_weight[191][69],
reservoir_weight[191][70],
reservoir_weight[191][71],
reservoir_weight[191][72],
reservoir_weight[191][73],
reservoir_weight[191][74],
reservoir_weight[191][75],
reservoir_weight[191][76],
reservoir_weight[191][77],
reservoir_weight[191][78],
reservoir_weight[191][79],
reservoir_weight[191][80],
reservoir_weight[191][81],
reservoir_weight[191][82],
reservoir_weight[191][83],
reservoir_weight[191][84],
reservoir_weight[191][85],
reservoir_weight[191][86],
reservoir_weight[191][87],
reservoir_weight[191][88],
reservoir_weight[191][89],
reservoir_weight[191][90],
reservoir_weight[191][91],
reservoir_weight[191][92],
reservoir_weight[191][93],
reservoir_weight[191][94],
reservoir_weight[191][95],
reservoir_weight[191][96],
reservoir_weight[191][97],
reservoir_weight[191][98],
reservoir_weight[191][99],
reservoir_weight[191][100],
reservoir_weight[191][101],
reservoir_weight[191][102],
reservoir_weight[191][103],
reservoir_weight[191][104],
reservoir_weight[191][105],
reservoir_weight[191][106],
reservoir_weight[191][107],
reservoir_weight[191][108],
reservoir_weight[191][109],
reservoir_weight[191][110],
reservoir_weight[191][111],
reservoir_weight[191][112],
reservoir_weight[191][113],
reservoir_weight[191][114],
reservoir_weight[191][115],
reservoir_weight[191][116],
reservoir_weight[191][117],
reservoir_weight[191][118],
reservoir_weight[191][119],
reservoir_weight[191][120],
reservoir_weight[191][121],
reservoir_weight[191][122],
reservoir_weight[191][123],
reservoir_weight[191][124],
reservoir_weight[191][125],
reservoir_weight[191][126],
reservoir_weight[191][127],
reservoir_weight[191][128],
reservoir_weight[191][129],
reservoir_weight[191][130],
reservoir_weight[191][131],
reservoir_weight[191][132],
reservoir_weight[191][133],
reservoir_weight[191][134],
reservoir_weight[191][135],
reservoir_weight[191][136],
reservoir_weight[191][137],
reservoir_weight[191][138],
reservoir_weight[191][139],
reservoir_weight[191][140],
reservoir_weight[191][141],
reservoir_weight[191][142],
reservoir_weight[191][143],
reservoir_weight[191][144],
reservoir_weight[191][145],
reservoir_weight[191][146],
reservoir_weight[191][147],
reservoir_weight[191][148],
reservoir_weight[191][149],
reservoir_weight[191][150],
reservoir_weight[191][151],
reservoir_weight[191][152],
reservoir_weight[191][153],
reservoir_weight[191][154],
reservoir_weight[191][155],
reservoir_weight[191][156],
reservoir_weight[191][157],
reservoir_weight[191][158],
reservoir_weight[191][159],
reservoir_weight[191][160],
reservoir_weight[191][161],
reservoir_weight[191][162],
reservoir_weight[191][163],
reservoir_weight[191][164],
reservoir_weight[191][165],
reservoir_weight[191][166],
reservoir_weight[191][167],
reservoir_weight[191][168],
reservoir_weight[191][169],
reservoir_weight[191][170],
reservoir_weight[191][171],
reservoir_weight[191][172],
reservoir_weight[191][173],
reservoir_weight[191][174],
reservoir_weight[191][175],
reservoir_weight[191][176],
reservoir_weight[191][177],
reservoir_weight[191][178],
reservoir_weight[191][179],
reservoir_weight[191][180],
reservoir_weight[191][181],
reservoir_weight[191][182],
reservoir_weight[191][183],
reservoir_weight[191][184],
reservoir_weight[191][185],
reservoir_weight[191][186],
reservoir_weight[191][187],
reservoir_weight[191][188],
reservoir_weight[191][189],
reservoir_weight[191][190],
reservoir_weight[191][191],
reservoir_weight[191][192],
reservoir_weight[191][193],
reservoir_weight[191][194],
reservoir_weight[191][195],
reservoir_weight[191][196],
reservoir_weight[191][197],
reservoir_weight[191][198],
reservoir_weight[191][199]
},
{reservoir_weight[192][0],
reservoir_weight[192][1],
reservoir_weight[192][2],
reservoir_weight[192][3],
reservoir_weight[192][4],
reservoir_weight[192][5],
reservoir_weight[192][6],
reservoir_weight[192][7],
reservoir_weight[192][8],
reservoir_weight[192][9],
reservoir_weight[192][10],
reservoir_weight[192][11],
reservoir_weight[192][12],
reservoir_weight[192][13],
reservoir_weight[192][14],
reservoir_weight[192][15],
reservoir_weight[192][16],
reservoir_weight[192][17],
reservoir_weight[192][18],
reservoir_weight[192][19],
reservoir_weight[192][20],
reservoir_weight[192][21],
reservoir_weight[192][22],
reservoir_weight[192][23],
reservoir_weight[192][24],
reservoir_weight[192][25],
reservoir_weight[192][26],
reservoir_weight[192][27],
reservoir_weight[192][28],
reservoir_weight[192][29],
reservoir_weight[192][30],
reservoir_weight[192][31],
reservoir_weight[192][32],
reservoir_weight[192][33],
reservoir_weight[192][34],
reservoir_weight[192][35],
reservoir_weight[192][36],
reservoir_weight[192][37],
reservoir_weight[192][38],
reservoir_weight[192][39],
reservoir_weight[192][40],
reservoir_weight[192][41],
reservoir_weight[192][42],
reservoir_weight[192][43],
reservoir_weight[192][44],
reservoir_weight[192][45],
reservoir_weight[192][46],
reservoir_weight[192][47],
reservoir_weight[192][48],
reservoir_weight[192][49],
reservoir_weight[192][50],
reservoir_weight[192][51],
reservoir_weight[192][52],
reservoir_weight[192][53],
reservoir_weight[192][54],
reservoir_weight[192][55],
reservoir_weight[192][56],
reservoir_weight[192][57],
reservoir_weight[192][58],
reservoir_weight[192][59],
reservoir_weight[192][60],
reservoir_weight[192][61],
reservoir_weight[192][62],
reservoir_weight[192][63],
reservoir_weight[192][64],
reservoir_weight[192][65],
reservoir_weight[192][66],
reservoir_weight[192][67],
reservoir_weight[192][68],
reservoir_weight[192][69],
reservoir_weight[192][70],
reservoir_weight[192][71],
reservoir_weight[192][72],
reservoir_weight[192][73],
reservoir_weight[192][74],
reservoir_weight[192][75],
reservoir_weight[192][76],
reservoir_weight[192][77],
reservoir_weight[192][78],
reservoir_weight[192][79],
reservoir_weight[192][80],
reservoir_weight[192][81],
reservoir_weight[192][82],
reservoir_weight[192][83],
reservoir_weight[192][84],
reservoir_weight[192][85],
reservoir_weight[192][86],
reservoir_weight[192][87],
reservoir_weight[192][88],
reservoir_weight[192][89],
reservoir_weight[192][90],
reservoir_weight[192][91],
reservoir_weight[192][92],
reservoir_weight[192][93],
reservoir_weight[192][94],
reservoir_weight[192][95],
reservoir_weight[192][96],
reservoir_weight[192][97],
reservoir_weight[192][98],
reservoir_weight[192][99],
reservoir_weight[192][100],
reservoir_weight[192][101],
reservoir_weight[192][102],
reservoir_weight[192][103],
reservoir_weight[192][104],
reservoir_weight[192][105],
reservoir_weight[192][106],
reservoir_weight[192][107],
reservoir_weight[192][108],
reservoir_weight[192][109],
reservoir_weight[192][110],
reservoir_weight[192][111],
reservoir_weight[192][112],
reservoir_weight[192][113],
reservoir_weight[192][114],
reservoir_weight[192][115],
reservoir_weight[192][116],
reservoir_weight[192][117],
reservoir_weight[192][118],
reservoir_weight[192][119],
reservoir_weight[192][120],
reservoir_weight[192][121],
reservoir_weight[192][122],
reservoir_weight[192][123],
reservoir_weight[192][124],
reservoir_weight[192][125],
reservoir_weight[192][126],
reservoir_weight[192][127],
reservoir_weight[192][128],
reservoir_weight[192][129],
reservoir_weight[192][130],
reservoir_weight[192][131],
reservoir_weight[192][132],
reservoir_weight[192][133],
reservoir_weight[192][134],
reservoir_weight[192][135],
reservoir_weight[192][136],
reservoir_weight[192][137],
reservoir_weight[192][138],
reservoir_weight[192][139],
reservoir_weight[192][140],
reservoir_weight[192][141],
reservoir_weight[192][142],
reservoir_weight[192][143],
reservoir_weight[192][144],
reservoir_weight[192][145],
reservoir_weight[192][146],
reservoir_weight[192][147],
reservoir_weight[192][148],
reservoir_weight[192][149],
reservoir_weight[192][150],
reservoir_weight[192][151],
reservoir_weight[192][152],
reservoir_weight[192][153],
reservoir_weight[192][154],
reservoir_weight[192][155],
reservoir_weight[192][156],
reservoir_weight[192][157],
reservoir_weight[192][158],
reservoir_weight[192][159],
reservoir_weight[192][160],
reservoir_weight[192][161],
reservoir_weight[192][162],
reservoir_weight[192][163],
reservoir_weight[192][164],
reservoir_weight[192][165],
reservoir_weight[192][166],
reservoir_weight[192][167],
reservoir_weight[192][168],
reservoir_weight[192][169],
reservoir_weight[192][170],
reservoir_weight[192][171],
reservoir_weight[192][172],
reservoir_weight[192][173],
reservoir_weight[192][174],
reservoir_weight[192][175],
reservoir_weight[192][176],
reservoir_weight[192][177],
reservoir_weight[192][178],
reservoir_weight[192][179],
reservoir_weight[192][180],
reservoir_weight[192][181],
reservoir_weight[192][182],
reservoir_weight[192][183],
reservoir_weight[192][184],
reservoir_weight[192][185],
reservoir_weight[192][186],
reservoir_weight[192][187],
reservoir_weight[192][188],
reservoir_weight[192][189],
reservoir_weight[192][190],
reservoir_weight[192][191],
reservoir_weight[192][192],
reservoir_weight[192][193],
reservoir_weight[192][194],
reservoir_weight[192][195],
reservoir_weight[192][196],
reservoir_weight[192][197],
reservoir_weight[192][198],
reservoir_weight[192][199]
},
{reservoir_weight[193][0],
reservoir_weight[193][1],
reservoir_weight[193][2],
reservoir_weight[193][3],
reservoir_weight[193][4],
reservoir_weight[193][5],
reservoir_weight[193][6],
reservoir_weight[193][7],
reservoir_weight[193][8],
reservoir_weight[193][9],
reservoir_weight[193][10],
reservoir_weight[193][11],
reservoir_weight[193][12],
reservoir_weight[193][13],
reservoir_weight[193][14],
reservoir_weight[193][15],
reservoir_weight[193][16],
reservoir_weight[193][17],
reservoir_weight[193][18],
reservoir_weight[193][19],
reservoir_weight[193][20],
reservoir_weight[193][21],
reservoir_weight[193][22],
reservoir_weight[193][23],
reservoir_weight[193][24],
reservoir_weight[193][25],
reservoir_weight[193][26],
reservoir_weight[193][27],
reservoir_weight[193][28],
reservoir_weight[193][29],
reservoir_weight[193][30],
reservoir_weight[193][31],
reservoir_weight[193][32],
reservoir_weight[193][33],
reservoir_weight[193][34],
reservoir_weight[193][35],
reservoir_weight[193][36],
reservoir_weight[193][37],
reservoir_weight[193][38],
reservoir_weight[193][39],
reservoir_weight[193][40],
reservoir_weight[193][41],
reservoir_weight[193][42],
reservoir_weight[193][43],
reservoir_weight[193][44],
reservoir_weight[193][45],
reservoir_weight[193][46],
reservoir_weight[193][47],
reservoir_weight[193][48],
reservoir_weight[193][49],
reservoir_weight[193][50],
reservoir_weight[193][51],
reservoir_weight[193][52],
reservoir_weight[193][53],
reservoir_weight[193][54],
reservoir_weight[193][55],
reservoir_weight[193][56],
reservoir_weight[193][57],
reservoir_weight[193][58],
reservoir_weight[193][59],
reservoir_weight[193][60],
reservoir_weight[193][61],
reservoir_weight[193][62],
reservoir_weight[193][63],
reservoir_weight[193][64],
reservoir_weight[193][65],
reservoir_weight[193][66],
reservoir_weight[193][67],
reservoir_weight[193][68],
reservoir_weight[193][69],
reservoir_weight[193][70],
reservoir_weight[193][71],
reservoir_weight[193][72],
reservoir_weight[193][73],
reservoir_weight[193][74],
reservoir_weight[193][75],
reservoir_weight[193][76],
reservoir_weight[193][77],
reservoir_weight[193][78],
reservoir_weight[193][79],
reservoir_weight[193][80],
reservoir_weight[193][81],
reservoir_weight[193][82],
reservoir_weight[193][83],
reservoir_weight[193][84],
reservoir_weight[193][85],
reservoir_weight[193][86],
reservoir_weight[193][87],
reservoir_weight[193][88],
reservoir_weight[193][89],
reservoir_weight[193][90],
reservoir_weight[193][91],
reservoir_weight[193][92],
reservoir_weight[193][93],
reservoir_weight[193][94],
reservoir_weight[193][95],
reservoir_weight[193][96],
reservoir_weight[193][97],
reservoir_weight[193][98],
reservoir_weight[193][99],
reservoir_weight[193][100],
reservoir_weight[193][101],
reservoir_weight[193][102],
reservoir_weight[193][103],
reservoir_weight[193][104],
reservoir_weight[193][105],
reservoir_weight[193][106],
reservoir_weight[193][107],
reservoir_weight[193][108],
reservoir_weight[193][109],
reservoir_weight[193][110],
reservoir_weight[193][111],
reservoir_weight[193][112],
reservoir_weight[193][113],
reservoir_weight[193][114],
reservoir_weight[193][115],
reservoir_weight[193][116],
reservoir_weight[193][117],
reservoir_weight[193][118],
reservoir_weight[193][119],
reservoir_weight[193][120],
reservoir_weight[193][121],
reservoir_weight[193][122],
reservoir_weight[193][123],
reservoir_weight[193][124],
reservoir_weight[193][125],
reservoir_weight[193][126],
reservoir_weight[193][127],
reservoir_weight[193][128],
reservoir_weight[193][129],
reservoir_weight[193][130],
reservoir_weight[193][131],
reservoir_weight[193][132],
reservoir_weight[193][133],
reservoir_weight[193][134],
reservoir_weight[193][135],
reservoir_weight[193][136],
reservoir_weight[193][137],
reservoir_weight[193][138],
reservoir_weight[193][139],
reservoir_weight[193][140],
reservoir_weight[193][141],
reservoir_weight[193][142],
reservoir_weight[193][143],
reservoir_weight[193][144],
reservoir_weight[193][145],
reservoir_weight[193][146],
reservoir_weight[193][147],
reservoir_weight[193][148],
reservoir_weight[193][149],
reservoir_weight[193][150],
reservoir_weight[193][151],
reservoir_weight[193][152],
reservoir_weight[193][153],
reservoir_weight[193][154],
reservoir_weight[193][155],
reservoir_weight[193][156],
reservoir_weight[193][157],
reservoir_weight[193][158],
reservoir_weight[193][159],
reservoir_weight[193][160],
reservoir_weight[193][161],
reservoir_weight[193][162],
reservoir_weight[193][163],
reservoir_weight[193][164],
reservoir_weight[193][165],
reservoir_weight[193][166],
reservoir_weight[193][167],
reservoir_weight[193][168],
reservoir_weight[193][169],
reservoir_weight[193][170],
reservoir_weight[193][171],
reservoir_weight[193][172],
reservoir_weight[193][173],
reservoir_weight[193][174],
reservoir_weight[193][175],
reservoir_weight[193][176],
reservoir_weight[193][177],
reservoir_weight[193][178],
reservoir_weight[193][179],
reservoir_weight[193][180],
reservoir_weight[193][181],
reservoir_weight[193][182],
reservoir_weight[193][183],
reservoir_weight[193][184],
reservoir_weight[193][185],
reservoir_weight[193][186],
reservoir_weight[193][187],
reservoir_weight[193][188],
reservoir_weight[193][189],
reservoir_weight[193][190],
reservoir_weight[193][191],
reservoir_weight[193][192],
reservoir_weight[193][193],
reservoir_weight[193][194],
reservoir_weight[193][195],
reservoir_weight[193][196],
reservoir_weight[193][197],
reservoir_weight[193][198],
reservoir_weight[193][199]
},
{reservoir_weight[194][0],
reservoir_weight[194][1],
reservoir_weight[194][2],
reservoir_weight[194][3],
reservoir_weight[194][4],
reservoir_weight[194][5],
reservoir_weight[194][6],
reservoir_weight[194][7],
reservoir_weight[194][8],
reservoir_weight[194][9],
reservoir_weight[194][10],
reservoir_weight[194][11],
reservoir_weight[194][12],
reservoir_weight[194][13],
reservoir_weight[194][14],
reservoir_weight[194][15],
reservoir_weight[194][16],
reservoir_weight[194][17],
reservoir_weight[194][18],
reservoir_weight[194][19],
reservoir_weight[194][20],
reservoir_weight[194][21],
reservoir_weight[194][22],
reservoir_weight[194][23],
reservoir_weight[194][24],
reservoir_weight[194][25],
reservoir_weight[194][26],
reservoir_weight[194][27],
reservoir_weight[194][28],
reservoir_weight[194][29],
reservoir_weight[194][30],
reservoir_weight[194][31],
reservoir_weight[194][32],
reservoir_weight[194][33],
reservoir_weight[194][34],
reservoir_weight[194][35],
reservoir_weight[194][36],
reservoir_weight[194][37],
reservoir_weight[194][38],
reservoir_weight[194][39],
reservoir_weight[194][40],
reservoir_weight[194][41],
reservoir_weight[194][42],
reservoir_weight[194][43],
reservoir_weight[194][44],
reservoir_weight[194][45],
reservoir_weight[194][46],
reservoir_weight[194][47],
reservoir_weight[194][48],
reservoir_weight[194][49],
reservoir_weight[194][50],
reservoir_weight[194][51],
reservoir_weight[194][52],
reservoir_weight[194][53],
reservoir_weight[194][54],
reservoir_weight[194][55],
reservoir_weight[194][56],
reservoir_weight[194][57],
reservoir_weight[194][58],
reservoir_weight[194][59],
reservoir_weight[194][60],
reservoir_weight[194][61],
reservoir_weight[194][62],
reservoir_weight[194][63],
reservoir_weight[194][64],
reservoir_weight[194][65],
reservoir_weight[194][66],
reservoir_weight[194][67],
reservoir_weight[194][68],
reservoir_weight[194][69],
reservoir_weight[194][70],
reservoir_weight[194][71],
reservoir_weight[194][72],
reservoir_weight[194][73],
reservoir_weight[194][74],
reservoir_weight[194][75],
reservoir_weight[194][76],
reservoir_weight[194][77],
reservoir_weight[194][78],
reservoir_weight[194][79],
reservoir_weight[194][80],
reservoir_weight[194][81],
reservoir_weight[194][82],
reservoir_weight[194][83],
reservoir_weight[194][84],
reservoir_weight[194][85],
reservoir_weight[194][86],
reservoir_weight[194][87],
reservoir_weight[194][88],
reservoir_weight[194][89],
reservoir_weight[194][90],
reservoir_weight[194][91],
reservoir_weight[194][92],
reservoir_weight[194][93],
reservoir_weight[194][94],
reservoir_weight[194][95],
reservoir_weight[194][96],
reservoir_weight[194][97],
reservoir_weight[194][98],
reservoir_weight[194][99],
reservoir_weight[194][100],
reservoir_weight[194][101],
reservoir_weight[194][102],
reservoir_weight[194][103],
reservoir_weight[194][104],
reservoir_weight[194][105],
reservoir_weight[194][106],
reservoir_weight[194][107],
reservoir_weight[194][108],
reservoir_weight[194][109],
reservoir_weight[194][110],
reservoir_weight[194][111],
reservoir_weight[194][112],
reservoir_weight[194][113],
reservoir_weight[194][114],
reservoir_weight[194][115],
reservoir_weight[194][116],
reservoir_weight[194][117],
reservoir_weight[194][118],
reservoir_weight[194][119],
reservoir_weight[194][120],
reservoir_weight[194][121],
reservoir_weight[194][122],
reservoir_weight[194][123],
reservoir_weight[194][124],
reservoir_weight[194][125],
reservoir_weight[194][126],
reservoir_weight[194][127],
reservoir_weight[194][128],
reservoir_weight[194][129],
reservoir_weight[194][130],
reservoir_weight[194][131],
reservoir_weight[194][132],
reservoir_weight[194][133],
reservoir_weight[194][134],
reservoir_weight[194][135],
reservoir_weight[194][136],
reservoir_weight[194][137],
reservoir_weight[194][138],
reservoir_weight[194][139],
reservoir_weight[194][140],
reservoir_weight[194][141],
reservoir_weight[194][142],
reservoir_weight[194][143],
reservoir_weight[194][144],
reservoir_weight[194][145],
reservoir_weight[194][146],
reservoir_weight[194][147],
reservoir_weight[194][148],
reservoir_weight[194][149],
reservoir_weight[194][150],
reservoir_weight[194][151],
reservoir_weight[194][152],
reservoir_weight[194][153],
reservoir_weight[194][154],
reservoir_weight[194][155],
reservoir_weight[194][156],
reservoir_weight[194][157],
reservoir_weight[194][158],
reservoir_weight[194][159],
reservoir_weight[194][160],
reservoir_weight[194][161],
reservoir_weight[194][162],
reservoir_weight[194][163],
reservoir_weight[194][164],
reservoir_weight[194][165],
reservoir_weight[194][166],
reservoir_weight[194][167],
reservoir_weight[194][168],
reservoir_weight[194][169],
reservoir_weight[194][170],
reservoir_weight[194][171],
reservoir_weight[194][172],
reservoir_weight[194][173],
reservoir_weight[194][174],
reservoir_weight[194][175],
reservoir_weight[194][176],
reservoir_weight[194][177],
reservoir_weight[194][178],
reservoir_weight[194][179],
reservoir_weight[194][180],
reservoir_weight[194][181],
reservoir_weight[194][182],
reservoir_weight[194][183],
reservoir_weight[194][184],
reservoir_weight[194][185],
reservoir_weight[194][186],
reservoir_weight[194][187],
reservoir_weight[194][188],
reservoir_weight[194][189],
reservoir_weight[194][190],
reservoir_weight[194][191],
reservoir_weight[194][192],
reservoir_weight[194][193],
reservoir_weight[194][194],
reservoir_weight[194][195],
reservoir_weight[194][196],
reservoir_weight[194][197],
reservoir_weight[194][198],
reservoir_weight[194][199]
},
{reservoir_weight[195][0],
reservoir_weight[195][1],
reservoir_weight[195][2],
reservoir_weight[195][3],
reservoir_weight[195][4],
reservoir_weight[195][5],
reservoir_weight[195][6],
reservoir_weight[195][7],
reservoir_weight[195][8],
reservoir_weight[195][9],
reservoir_weight[195][10],
reservoir_weight[195][11],
reservoir_weight[195][12],
reservoir_weight[195][13],
reservoir_weight[195][14],
reservoir_weight[195][15],
reservoir_weight[195][16],
reservoir_weight[195][17],
reservoir_weight[195][18],
reservoir_weight[195][19],
reservoir_weight[195][20],
reservoir_weight[195][21],
reservoir_weight[195][22],
reservoir_weight[195][23],
reservoir_weight[195][24],
reservoir_weight[195][25],
reservoir_weight[195][26],
reservoir_weight[195][27],
reservoir_weight[195][28],
reservoir_weight[195][29],
reservoir_weight[195][30],
reservoir_weight[195][31],
reservoir_weight[195][32],
reservoir_weight[195][33],
reservoir_weight[195][34],
reservoir_weight[195][35],
reservoir_weight[195][36],
reservoir_weight[195][37],
reservoir_weight[195][38],
reservoir_weight[195][39],
reservoir_weight[195][40],
reservoir_weight[195][41],
reservoir_weight[195][42],
reservoir_weight[195][43],
reservoir_weight[195][44],
reservoir_weight[195][45],
reservoir_weight[195][46],
reservoir_weight[195][47],
reservoir_weight[195][48],
reservoir_weight[195][49],
reservoir_weight[195][50],
reservoir_weight[195][51],
reservoir_weight[195][52],
reservoir_weight[195][53],
reservoir_weight[195][54],
reservoir_weight[195][55],
reservoir_weight[195][56],
reservoir_weight[195][57],
reservoir_weight[195][58],
reservoir_weight[195][59],
reservoir_weight[195][60],
reservoir_weight[195][61],
reservoir_weight[195][62],
reservoir_weight[195][63],
reservoir_weight[195][64],
reservoir_weight[195][65],
reservoir_weight[195][66],
reservoir_weight[195][67],
reservoir_weight[195][68],
reservoir_weight[195][69],
reservoir_weight[195][70],
reservoir_weight[195][71],
reservoir_weight[195][72],
reservoir_weight[195][73],
reservoir_weight[195][74],
reservoir_weight[195][75],
reservoir_weight[195][76],
reservoir_weight[195][77],
reservoir_weight[195][78],
reservoir_weight[195][79],
reservoir_weight[195][80],
reservoir_weight[195][81],
reservoir_weight[195][82],
reservoir_weight[195][83],
reservoir_weight[195][84],
reservoir_weight[195][85],
reservoir_weight[195][86],
reservoir_weight[195][87],
reservoir_weight[195][88],
reservoir_weight[195][89],
reservoir_weight[195][90],
reservoir_weight[195][91],
reservoir_weight[195][92],
reservoir_weight[195][93],
reservoir_weight[195][94],
reservoir_weight[195][95],
reservoir_weight[195][96],
reservoir_weight[195][97],
reservoir_weight[195][98],
reservoir_weight[195][99],
reservoir_weight[195][100],
reservoir_weight[195][101],
reservoir_weight[195][102],
reservoir_weight[195][103],
reservoir_weight[195][104],
reservoir_weight[195][105],
reservoir_weight[195][106],
reservoir_weight[195][107],
reservoir_weight[195][108],
reservoir_weight[195][109],
reservoir_weight[195][110],
reservoir_weight[195][111],
reservoir_weight[195][112],
reservoir_weight[195][113],
reservoir_weight[195][114],
reservoir_weight[195][115],
reservoir_weight[195][116],
reservoir_weight[195][117],
reservoir_weight[195][118],
reservoir_weight[195][119],
reservoir_weight[195][120],
reservoir_weight[195][121],
reservoir_weight[195][122],
reservoir_weight[195][123],
reservoir_weight[195][124],
reservoir_weight[195][125],
reservoir_weight[195][126],
reservoir_weight[195][127],
reservoir_weight[195][128],
reservoir_weight[195][129],
reservoir_weight[195][130],
reservoir_weight[195][131],
reservoir_weight[195][132],
reservoir_weight[195][133],
reservoir_weight[195][134],
reservoir_weight[195][135],
reservoir_weight[195][136],
reservoir_weight[195][137],
reservoir_weight[195][138],
reservoir_weight[195][139],
reservoir_weight[195][140],
reservoir_weight[195][141],
reservoir_weight[195][142],
reservoir_weight[195][143],
reservoir_weight[195][144],
reservoir_weight[195][145],
reservoir_weight[195][146],
reservoir_weight[195][147],
reservoir_weight[195][148],
reservoir_weight[195][149],
reservoir_weight[195][150],
reservoir_weight[195][151],
reservoir_weight[195][152],
reservoir_weight[195][153],
reservoir_weight[195][154],
reservoir_weight[195][155],
reservoir_weight[195][156],
reservoir_weight[195][157],
reservoir_weight[195][158],
reservoir_weight[195][159],
reservoir_weight[195][160],
reservoir_weight[195][161],
reservoir_weight[195][162],
reservoir_weight[195][163],
reservoir_weight[195][164],
reservoir_weight[195][165],
reservoir_weight[195][166],
reservoir_weight[195][167],
reservoir_weight[195][168],
reservoir_weight[195][169],
reservoir_weight[195][170],
reservoir_weight[195][171],
reservoir_weight[195][172],
reservoir_weight[195][173],
reservoir_weight[195][174],
reservoir_weight[195][175],
reservoir_weight[195][176],
reservoir_weight[195][177],
reservoir_weight[195][178],
reservoir_weight[195][179],
reservoir_weight[195][180],
reservoir_weight[195][181],
reservoir_weight[195][182],
reservoir_weight[195][183],
reservoir_weight[195][184],
reservoir_weight[195][185],
reservoir_weight[195][186],
reservoir_weight[195][187],
reservoir_weight[195][188],
reservoir_weight[195][189],
reservoir_weight[195][190],
reservoir_weight[195][191],
reservoir_weight[195][192],
reservoir_weight[195][193],
reservoir_weight[195][194],
reservoir_weight[195][195],
reservoir_weight[195][196],
reservoir_weight[195][197],
reservoir_weight[195][198],
reservoir_weight[195][199]
},
{reservoir_weight[196][0],
reservoir_weight[196][1],
reservoir_weight[196][2],
reservoir_weight[196][3],
reservoir_weight[196][4],
reservoir_weight[196][5],
reservoir_weight[196][6],
reservoir_weight[196][7],
reservoir_weight[196][8],
reservoir_weight[196][9],
reservoir_weight[196][10],
reservoir_weight[196][11],
reservoir_weight[196][12],
reservoir_weight[196][13],
reservoir_weight[196][14],
reservoir_weight[196][15],
reservoir_weight[196][16],
reservoir_weight[196][17],
reservoir_weight[196][18],
reservoir_weight[196][19],
reservoir_weight[196][20],
reservoir_weight[196][21],
reservoir_weight[196][22],
reservoir_weight[196][23],
reservoir_weight[196][24],
reservoir_weight[196][25],
reservoir_weight[196][26],
reservoir_weight[196][27],
reservoir_weight[196][28],
reservoir_weight[196][29],
reservoir_weight[196][30],
reservoir_weight[196][31],
reservoir_weight[196][32],
reservoir_weight[196][33],
reservoir_weight[196][34],
reservoir_weight[196][35],
reservoir_weight[196][36],
reservoir_weight[196][37],
reservoir_weight[196][38],
reservoir_weight[196][39],
reservoir_weight[196][40],
reservoir_weight[196][41],
reservoir_weight[196][42],
reservoir_weight[196][43],
reservoir_weight[196][44],
reservoir_weight[196][45],
reservoir_weight[196][46],
reservoir_weight[196][47],
reservoir_weight[196][48],
reservoir_weight[196][49],
reservoir_weight[196][50],
reservoir_weight[196][51],
reservoir_weight[196][52],
reservoir_weight[196][53],
reservoir_weight[196][54],
reservoir_weight[196][55],
reservoir_weight[196][56],
reservoir_weight[196][57],
reservoir_weight[196][58],
reservoir_weight[196][59],
reservoir_weight[196][60],
reservoir_weight[196][61],
reservoir_weight[196][62],
reservoir_weight[196][63],
reservoir_weight[196][64],
reservoir_weight[196][65],
reservoir_weight[196][66],
reservoir_weight[196][67],
reservoir_weight[196][68],
reservoir_weight[196][69],
reservoir_weight[196][70],
reservoir_weight[196][71],
reservoir_weight[196][72],
reservoir_weight[196][73],
reservoir_weight[196][74],
reservoir_weight[196][75],
reservoir_weight[196][76],
reservoir_weight[196][77],
reservoir_weight[196][78],
reservoir_weight[196][79],
reservoir_weight[196][80],
reservoir_weight[196][81],
reservoir_weight[196][82],
reservoir_weight[196][83],
reservoir_weight[196][84],
reservoir_weight[196][85],
reservoir_weight[196][86],
reservoir_weight[196][87],
reservoir_weight[196][88],
reservoir_weight[196][89],
reservoir_weight[196][90],
reservoir_weight[196][91],
reservoir_weight[196][92],
reservoir_weight[196][93],
reservoir_weight[196][94],
reservoir_weight[196][95],
reservoir_weight[196][96],
reservoir_weight[196][97],
reservoir_weight[196][98],
reservoir_weight[196][99],
reservoir_weight[196][100],
reservoir_weight[196][101],
reservoir_weight[196][102],
reservoir_weight[196][103],
reservoir_weight[196][104],
reservoir_weight[196][105],
reservoir_weight[196][106],
reservoir_weight[196][107],
reservoir_weight[196][108],
reservoir_weight[196][109],
reservoir_weight[196][110],
reservoir_weight[196][111],
reservoir_weight[196][112],
reservoir_weight[196][113],
reservoir_weight[196][114],
reservoir_weight[196][115],
reservoir_weight[196][116],
reservoir_weight[196][117],
reservoir_weight[196][118],
reservoir_weight[196][119],
reservoir_weight[196][120],
reservoir_weight[196][121],
reservoir_weight[196][122],
reservoir_weight[196][123],
reservoir_weight[196][124],
reservoir_weight[196][125],
reservoir_weight[196][126],
reservoir_weight[196][127],
reservoir_weight[196][128],
reservoir_weight[196][129],
reservoir_weight[196][130],
reservoir_weight[196][131],
reservoir_weight[196][132],
reservoir_weight[196][133],
reservoir_weight[196][134],
reservoir_weight[196][135],
reservoir_weight[196][136],
reservoir_weight[196][137],
reservoir_weight[196][138],
reservoir_weight[196][139],
reservoir_weight[196][140],
reservoir_weight[196][141],
reservoir_weight[196][142],
reservoir_weight[196][143],
reservoir_weight[196][144],
reservoir_weight[196][145],
reservoir_weight[196][146],
reservoir_weight[196][147],
reservoir_weight[196][148],
reservoir_weight[196][149],
reservoir_weight[196][150],
reservoir_weight[196][151],
reservoir_weight[196][152],
reservoir_weight[196][153],
reservoir_weight[196][154],
reservoir_weight[196][155],
reservoir_weight[196][156],
reservoir_weight[196][157],
reservoir_weight[196][158],
reservoir_weight[196][159],
reservoir_weight[196][160],
reservoir_weight[196][161],
reservoir_weight[196][162],
reservoir_weight[196][163],
reservoir_weight[196][164],
reservoir_weight[196][165],
reservoir_weight[196][166],
reservoir_weight[196][167],
reservoir_weight[196][168],
reservoir_weight[196][169],
reservoir_weight[196][170],
reservoir_weight[196][171],
reservoir_weight[196][172],
reservoir_weight[196][173],
reservoir_weight[196][174],
reservoir_weight[196][175],
reservoir_weight[196][176],
reservoir_weight[196][177],
reservoir_weight[196][178],
reservoir_weight[196][179],
reservoir_weight[196][180],
reservoir_weight[196][181],
reservoir_weight[196][182],
reservoir_weight[196][183],
reservoir_weight[196][184],
reservoir_weight[196][185],
reservoir_weight[196][186],
reservoir_weight[196][187],
reservoir_weight[196][188],
reservoir_weight[196][189],
reservoir_weight[196][190],
reservoir_weight[196][191],
reservoir_weight[196][192],
reservoir_weight[196][193],
reservoir_weight[196][194],
reservoir_weight[196][195],
reservoir_weight[196][196],
reservoir_weight[196][197],
reservoir_weight[196][198],
reservoir_weight[196][199]
},
{reservoir_weight[197][0],
reservoir_weight[197][1],
reservoir_weight[197][2],
reservoir_weight[197][3],
reservoir_weight[197][4],
reservoir_weight[197][5],
reservoir_weight[197][6],
reservoir_weight[197][7],
reservoir_weight[197][8],
reservoir_weight[197][9],
reservoir_weight[197][10],
reservoir_weight[197][11],
reservoir_weight[197][12],
reservoir_weight[197][13],
reservoir_weight[197][14],
reservoir_weight[197][15],
reservoir_weight[197][16],
reservoir_weight[197][17],
reservoir_weight[197][18],
reservoir_weight[197][19],
reservoir_weight[197][20],
reservoir_weight[197][21],
reservoir_weight[197][22],
reservoir_weight[197][23],
reservoir_weight[197][24],
reservoir_weight[197][25],
reservoir_weight[197][26],
reservoir_weight[197][27],
reservoir_weight[197][28],
reservoir_weight[197][29],
reservoir_weight[197][30],
reservoir_weight[197][31],
reservoir_weight[197][32],
reservoir_weight[197][33],
reservoir_weight[197][34],
reservoir_weight[197][35],
reservoir_weight[197][36],
reservoir_weight[197][37],
reservoir_weight[197][38],
reservoir_weight[197][39],
reservoir_weight[197][40],
reservoir_weight[197][41],
reservoir_weight[197][42],
reservoir_weight[197][43],
reservoir_weight[197][44],
reservoir_weight[197][45],
reservoir_weight[197][46],
reservoir_weight[197][47],
reservoir_weight[197][48],
reservoir_weight[197][49],
reservoir_weight[197][50],
reservoir_weight[197][51],
reservoir_weight[197][52],
reservoir_weight[197][53],
reservoir_weight[197][54],
reservoir_weight[197][55],
reservoir_weight[197][56],
reservoir_weight[197][57],
reservoir_weight[197][58],
reservoir_weight[197][59],
reservoir_weight[197][60],
reservoir_weight[197][61],
reservoir_weight[197][62],
reservoir_weight[197][63],
reservoir_weight[197][64],
reservoir_weight[197][65],
reservoir_weight[197][66],
reservoir_weight[197][67],
reservoir_weight[197][68],
reservoir_weight[197][69],
reservoir_weight[197][70],
reservoir_weight[197][71],
reservoir_weight[197][72],
reservoir_weight[197][73],
reservoir_weight[197][74],
reservoir_weight[197][75],
reservoir_weight[197][76],
reservoir_weight[197][77],
reservoir_weight[197][78],
reservoir_weight[197][79],
reservoir_weight[197][80],
reservoir_weight[197][81],
reservoir_weight[197][82],
reservoir_weight[197][83],
reservoir_weight[197][84],
reservoir_weight[197][85],
reservoir_weight[197][86],
reservoir_weight[197][87],
reservoir_weight[197][88],
reservoir_weight[197][89],
reservoir_weight[197][90],
reservoir_weight[197][91],
reservoir_weight[197][92],
reservoir_weight[197][93],
reservoir_weight[197][94],
reservoir_weight[197][95],
reservoir_weight[197][96],
reservoir_weight[197][97],
reservoir_weight[197][98],
reservoir_weight[197][99],
reservoir_weight[197][100],
reservoir_weight[197][101],
reservoir_weight[197][102],
reservoir_weight[197][103],
reservoir_weight[197][104],
reservoir_weight[197][105],
reservoir_weight[197][106],
reservoir_weight[197][107],
reservoir_weight[197][108],
reservoir_weight[197][109],
reservoir_weight[197][110],
reservoir_weight[197][111],
reservoir_weight[197][112],
reservoir_weight[197][113],
reservoir_weight[197][114],
reservoir_weight[197][115],
reservoir_weight[197][116],
reservoir_weight[197][117],
reservoir_weight[197][118],
reservoir_weight[197][119],
reservoir_weight[197][120],
reservoir_weight[197][121],
reservoir_weight[197][122],
reservoir_weight[197][123],
reservoir_weight[197][124],
reservoir_weight[197][125],
reservoir_weight[197][126],
reservoir_weight[197][127],
reservoir_weight[197][128],
reservoir_weight[197][129],
reservoir_weight[197][130],
reservoir_weight[197][131],
reservoir_weight[197][132],
reservoir_weight[197][133],
reservoir_weight[197][134],
reservoir_weight[197][135],
reservoir_weight[197][136],
reservoir_weight[197][137],
reservoir_weight[197][138],
reservoir_weight[197][139],
reservoir_weight[197][140],
reservoir_weight[197][141],
reservoir_weight[197][142],
reservoir_weight[197][143],
reservoir_weight[197][144],
reservoir_weight[197][145],
reservoir_weight[197][146],
reservoir_weight[197][147],
reservoir_weight[197][148],
reservoir_weight[197][149],
reservoir_weight[197][150],
reservoir_weight[197][151],
reservoir_weight[197][152],
reservoir_weight[197][153],
reservoir_weight[197][154],
reservoir_weight[197][155],
reservoir_weight[197][156],
reservoir_weight[197][157],
reservoir_weight[197][158],
reservoir_weight[197][159],
reservoir_weight[197][160],
reservoir_weight[197][161],
reservoir_weight[197][162],
reservoir_weight[197][163],
reservoir_weight[197][164],
reservoir_weight[197][165],
reservoir_weight[197][166],
reservoir_weight[197][167],
reservoir_weight[197][168],
reservoir_weight[197][169],
reservoir_weight[197][170],
reservoir_weight[197][171],
reservoir_weight[197][172],
reservoir_weight[197][173],
reservoir_weight[197][174],
reservoir_weight[197][175],
reservoir_weight[197][176],
reservoir_weight[197][177],
reservoir_weight[197][178],
reservoir_weight[197][179],
reservoir_weight[197][180],
reservoir_weight[197][181],
reservoir_weight[197][182],
reservoir_weight[197][183],
reservoir_weight[197][184],
reservoir_weight[197][185],
reservoir_weight[197][186],
reservoir_weight[197][187],
reservoir_weight[197][188],
reservoir_weight[197][189],
reservoir_weight[197][190],
reservoir_weight[197][191],
reservoir_weight[197][192],
reservoir_weight[197][193],
reservoir_weight[197][194],
reservoir_weight[197][195],
reservoir_weight[197][196],
reservoir_weight[197][197],
reservoir_weight[197][198],
reservoir_weight[197][199]
},
{reservoir_weight[198][0],
reservoir_weight[198][1],
reservoir_weight[198][2],
reservoir_weight[198][3],
reservoir_weight[198][4],
reservoir_weight[198][5],
reservoir_weight[198][6],
reservoir_weight[198][7],
reservoir_weight[198][8],
reservoir_weight[198][9],
reservoir_weight[198][10],
reservoir_weight[198][11],
reservoir_weight[198][12],
reservoir_weight[198][13],
reservoir_weight[198][14],
reservoir_weight[198][15],
reservoir_weight[198][16],
reservoir_weight[198][17],
reservoir_weight[198][18],
reservoir_weight[198][19],
reservoir_weight[198][20],
reservoir_weight[198][21],
reservoir_weight[198][22],
reservoir_weight[198][23],
reservoir_weight[198][24],
reservoir_weight[198][25],
reservoir_weight[198][26],
reservoir_weight[198][27],
reservoir_weight[198][28],
reservoir_weight[198][29],
reservoir_weight[198][30],
reservoir_weight[198][31],
reservoir_weight[198][32],
reservoir_weight[198][33],
reservoir_weight[198][34],
reservoir_weight[198][35],
reservoir_weight[198][36],
reservoir_weight[198][37],
reservoir_weight[198][38],
reservoir_weight[198][39],
reservoir_weight[198][40],
reservoir_weight[198][41],
reservoir_weight[198][42],
reservoir_weight[198][43],
reservoir_weight[198][44],
reservoir_weight[198][45],
reservoir_weight[198][46],
reservoir_weight[198][47],
reservoir_weight[198][48],
reservoir_weight[198][49],
reservoir_weight[198][50],
reservoir_weight[198][51],
reservoir_weight[198][52],
reservoir_weight[198][53],
reservoir_weight[198][54],
reservoir_weight[198][55],
reservoir_weight[198][56],
reservoir_weight[198][57],
reservoir_weight[198][58],
reservoir_weight[198][59],
reservoir_weight[198][60],
reservoir_weight[198][61],
reservoir_weight[198][62],
reservoir_weight[198][63],
reservoir_weight[198][64],
reservoir_weight[198][65],
reservoir_weight[198][66],
reservoir_weight[198][67],
reservoir_weight[198][68],
reservoir_weight[198][69],
reservoir_weight[198][70],
reservoir_weight[198][71],
reservoir_weight[198][72],
reservoir_weight[198][73],
reservoir_weight[198][74],
reservoir_weight[198][75],
reservoir_weight[198][76],
reservoir_weight[198][77],
reservoir_weight[198][78],
reservoir_weight[198][79],
reservoir_weight[198][80],
reservoir_weight[198][81],
reservoir_weight[198][82],
reservoir_weight[198][83],
reservoir_weight[198][84],
reservoir_weight[198][85],
reservoir_weight[198][86],
reservoir_weight[198][87],
reservoir_weight[198][88],
reservoir_weight[198][89],
reservoir_weight[198][90],
reservoir_weight[198][91],
reservoir_weight[198][92],
reservoir_weight[198][93],
reservoir_weight[198][94],
reservoir_weight[198][95],
reservoir_weight[198][96],
reservoir_weight[198][97],
reservoir_weight[198][98],
reservoir_weight[198][99],
reservoir_weight[198][100],
reservoir_weight[198][101],
reservoir_weight[198][102],
reservoir_weight[198][103],
reservoir_weight[198][104],
reservoir_weight[198][105],
reservoir_weight[198][106],
reservoir_weight[198][107],
reservoir_weight[198][108],
reservoir_weight[198][109],
reservoir_weight[198][110],
reservoir_weight[198][111],
reservoir_weight[198][112],
reservoir_weight[198][113],
reservoir_weight[198][114],
reservoir_weight[198][115],
reservoir_weight[198][116],
reservoir_weight[198][117],
reservoir_weight[198][118],
reservoir_weight[198][119],
reservoir_weight[198][120],
reservoir_weight[198][121],
reservoir_weight[198][122],
reservoir_weight[198][123],
reservoir_weight[198][124],
reservoir_weight[198][125],
reservoir_weight[198][126],
reservoir_weight[198][127],
reservoir_weight[198][128],
reservoir_weight[198][129],
reservoir_weight[198][130],
reservoir_weight[198][131],
reservoir_weight[198][132],
reservoir_weight[198][133],
reservoir_weight[198][134],
reservoir_weight[198][135],
reservoir_weight[198][136],
reservoir_weight[198][137],
reservoir_weight[198][138],
reservoir_weight[198][139],
reservoir_weight[198][140],
reservoir_weight[198][141],
reservoir_weight[198][142],
reservoir_weight[198][143],
reservoir_weight[198][144],
reservoir_weight[198][145],
reservoir_weight[198][146],
reservoir_weight[198][147],
reservoir_weight[198][148],
reservoir_weight[198][149],
reservoir_weight[198][150],
reservoir_weight[198][151],
reservoir_weight[198][152],
reservoir_weight[198][153],
reservoir_weight[198][154],
reservoir_weight[198][155],
reservoir_weight[198][156],
reservoir_weight[198][157],
reservoir_weight[198][158],
reservoir_weight[198][159],
reservoir_weight[198][160],
reservoir_weight[198][161],
reservoir_weight[198][162],
reservoir_weight[198][163],
reservoir_weight[198][164],
reservoir_weight[198][165],
reservoir_weight[198][166],
reservoir_weight[198][167],
reservoir_weight[198][168],
reservoir_weight[198][169],
reservoir_weight[198][170],
reservoir_weight[198][171],
reservoir_weight[198][172],
reservoir_weight[198][173],
reservoir_weight[198][174],
reservoir_weight[198][175],
reservoir_weight[198][176],
reservoir_weight[198][177],
reservoir_weight[198][178],
reservoir_weight[198][179],
reservoir_weight[198][180],
reservoir_weight[198][181],
reservoir_weight[198][182],
reservoir_weight[198][183],
reservoir_weight[198][184],
reservoir_weight[198][185],
reservoir_weight[198][186],
reservoir_weight[198][187],
reservoir_weight[198][188],
reservoir_weight[198][189],
reservoir_weight[198][190],
reservoir_weight[198][191],
reservoir_weight[198][192],
reservoir_weight[198][193],
reservoir_weight[198][194],
reservoir_weight[198][195],
reservoir_weight[198][196],
reservoir_weight[198][197],
reservoir_weight[198][198],
reservoir_weight[198][199]
},
{reservoir_weight[199][0],
reservoir_weight[199][1],
reservoir_weight[199][2],
reservoir_weight[199][3],
reservoir_weight[199][4],
reservoir_weight[199][5],
reservoir_weight[199][6],
reservoir_weight[199][7],
reservoir_weight[199][8],
reservoir_weight[199][9],
reservoir_weight[199][10],
reservoir_weight[199][11],
reservoir_weight[199][12],
reservoir_weight[199][13],
reservoir_weight[199][14],
reservoir_weight[199][15],
reservoir_weight[199][16],
reservoir_weight[199][17],
reservoir_weight[199][18],
reservoir_weight[199][19],
reservoir_weight[199][20],
reservoir_weight[199][21],
reservoir_weight[199][22],
reservoir_weight[199][23],
reservoir_weight[199][24],
reservoir_weight[199][25],
reservoir_weight[199][26],
reservoir_weight[199][27],
reservoir_weight[199][28],
reservoir_weight[199][29],
reservoir_weight[199][30],
reservoir_weight[199][31],
reservoir_weight[199][32],
reservoir_weight[199][33],
reservoir_weight[199][34],
reservoir_weight[199][35],
reservoir_weight[199][36],
reservoir_weight[199][37],
reservoir_weight[199][38],
reservoir_weight[199][39],
reservoir_weight[199][40],
reservoir_weight[199][41],
reservoir_weight[199][42],
reservoir_weight[199][43],
reservoir_weight[199][44],
reservoir_weight[199][45],
reservoir_weight[199][46],
reservoir_weight[199][47],
reservoir_weight[199][48],
reservoir_weight[199][49],
reservoir_weight[199][50],
reservoir_weight[199][51],
reservoir_weight[199][52],
reservoir_weight[199][53],
reservoir_weight[199][54],
reservoir_weight[199][55],
reservoir_weight[199][56],
reservoir_weight[199][57],
reservoir_weight[199][58],
reservoir_weight[199][59],
reservoir_weight[199][60],
reservoir_weight[199][61],
reservoir_weight[199][62],
reservoir_weight[199][63],
reservoir_weight[199][64],
reservoir_weight[199][65],
reservoir_weight[199][66],
reservoir_weight[199][67],
reservoir_weight[199][68],
reservoir_weight[199][69],
reservoir_weight[199][70],
reservoir_weight[199][71],
reservoir_weight[199][72],
reservoir_weight[199][73],
reservoir_weight[199][74],
reservoir_weight[199][75],
reservoir_weight[199][76],
reservoir_weight[199][77],
reservoir_weight[199][78],
reservoir_weight[199][79],
reservoir_weight[199][80],
reservoir_weight[199][81],
reservoir_weight[199][82],
reservoir_weight[199][83],
reservoir_weight[199][84],
reservoir_weight[199][85],
reservoir_weight[199][86],
reservoir_weight[199][87],
reservoir_weight[199][88],
reservoir_weight[199][89],
reservoir_weight[199][90],
reservoir_weight[199][91],
reservoir_weight[199][92],
reservoir_weight[199][93],
reservoir_weight[199][94],
reservoir_weight[199][95],
reservoir_weight[199][96],
reservoir_weight[199][97],
reservoir_weight[199][98],
reservoir_weight[199][99],
reservoir_weight[199][100],
reservoir_weight[199][101],
reservoir_weight[199][102],
reservoir_weight[199][103],
reservoir_weight[199][104],
reservoir_weight[199][105],
reservoir_weight[199][106],
reservoir_weight[199][107],
reservoir_weight[199][108],
reservoir_weight[199][109],
reservoir_weight[199][110],
reservoir_weight[199][111],
reservoir_weight[199][112],
reservoir_weight[199][113],
reservoir_weight[199][114],
reservoir_weight[199][115],
reservoir_weight[199][116],
reservoir_weight[199][117],
reservoir_weight[199][118],
reservoir_weight[199][119],
reservoir_weight[199][120],
reservoir_weight[199][121],
reservoir_weight[199][122],
reservoir_weight[199][123],
reservoir_weight[199][124],
reservoir_weight[199][125],
reservoir_weight[199][126],
reservoir_weight[199][127],
reservoir_weight[199][128],
reservoir_weight[199][129],
reservoir_weight[199][130],
reservoir_weight[199][131],
reservoir_weight[199][132],
reservoir_weight[199][133],
reservoir_weight[199][134],
reservoir_weight[199][135],
reservoir_weight[199][136],
reservoir_weight[199][137],
reservoir_weight[199][138],
reservoir_weight[199][139],
reservoir_weight[199][140],
reservoir_weight[199][141],
reservoir_weight[199][142],
reservoir_weight[199][143],
reservoir_weight[199][144],
reservoir_weight[199][145],
reservoir_weight[199][146],
reservoir_weight[199][147],
reservoir_weight[199][148],
reservoir_weight[199][149],
reservoir_weight[199][150],
reservoir_weight[199][151],
reservoir_weight[199][152],
reservoir_weight[199][153],
reservoir_weight[199][154],
reservoir_weight[199][155],
reservoir_weight[199][156],
reservoir_weight[199][157],
reservoir_weight[199][158],
reservoir_weight[199][159],
reservoir_weight[199][160],
reservoir_weight[199][161],
reservoir_weight[199][162],
reservoir_weight[199][163],
reservoir_weight[199][164],
reservoir_weight[199][165],
reservoir_weight[199][166],
reservoir_weight[199][167],
reservoir_weight[199][168],
reservoir_weight[199][169],
reservoir_weight[199][170],
reservoir_weight[199][171],
reservoir_weight[199][172],
reservoir_weight[199][173],
reservoir_weight[199][174],
reservoir_weight[199][175],
reservoir_weight[199][176],
reservoir_weight[199][177],
reservoir_weight[199][178],
reservoir_weight[199][179],
reservoir_weight[199][180],
reservoir_weight[199][181],
reservoir_weight[199][182],
reservoir_weight[199][183],
reservoir_weight[199][184],
reservoir_weight[199][185],
reservoir_weight[199][186],
reservoir_weight[199][187],
reservoir_weight[199][188],
reservoir_weight[199][189],
reservoir_weight[199][190],
reservoir_weight[199][191],
reservoir_weight[199][192],
reservoir_weight[199][193],
reservoir_weight[199][194],
reservoir_weight[199][195],
reservoir_weight[199][196],
reservoir_weight[199][197],
reservoir_weight[199][198],
reservoir_weight[199][199]
}
} = {
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
-8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd33,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd70,
-8'sd1,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd54,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
-8'sd13,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
-8'sd26,
-8'sd5,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd60,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd58,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd24,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
-8'sd80,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
-8'sd25,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd31,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
-8'sd47,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0
},
{8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
-8'sd13,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd73,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
-8'sd5,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0
},
{8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd70,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0,
8'sd0,
-8'sd11,
8'sd5,
8'sd68,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd57,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd42,
8'sd0,
-8'sd11,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd48,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd81,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
-8'sd62,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd29,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
-8'sd24,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
-8'sd9,
8'sd0,
8'sd22,
8'sd0,
8'sd7,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd69,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd70,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
-8'sd17,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
-8'sd45,
8'sd0,
-8'sd27,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd19,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
-8'sd64,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd58,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd79,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd75,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd61,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
-8'sd35,
8'sd5,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
-8'sd52,
8'sd0,
8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd42,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
-8'sd14,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd66,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
-8'sd24,
8'sd21,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd62,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd63,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
-8'sd31,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd45,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
-8'sd5,
8'sd0,
8'sd0,
-8'sd8,
8'sd5,
8'sd0,
8'sd4,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd59,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd49,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
-8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
-8'sd71,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
-8'sd11,
8'sd0,
8'sd27,
8'sd17,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd56,
8'sd0,
8'sd11,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd49,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd81,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd46,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd51,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd60,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
-8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd23,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd54,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd91,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd64,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
-8'sd54,
-8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd11,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd91,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd71,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd10,
8'sd67,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd45,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd89,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd65,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd0,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd57,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43
},
{8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd58,
8'sd0,
-8'sd34,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd73,
8'sd0,
-8'sd3,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd44,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd32,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd71,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
-8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd74,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
-8'sd19,
8'sd0,
-8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
-8'sd51,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd56,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd15,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd43,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd13,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd74,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd71,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd65,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
-8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd82,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd34,
8'sd16,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd67,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd39,
8'sd1,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd52,
8'sd0,
8'sd0,
-8'sd18,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd58,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd25,
8'sd61,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
-8'sd2,
8'sd10,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd66,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd77,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd52,
-8'sd8,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd56,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd71,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd80,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
-8'sd18,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd65,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd35,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd18,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd27,
-8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
-8'sd73,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd64,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{-8'sd79,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd23,
8'sd0,
8'sd0,
-8'sd46,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd42
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd63,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd74,
8'sd0,
-8'sd35,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd71,
8'sd68,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd54,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
-8'sd5,
-8'sd4,
8'sd0,
8'sd0,
-8'sd59,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd33,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
-8'sd14,
8'sd10,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
-8'sd31,
-8'sd10,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd88,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd49,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
-8'sd49,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
-8'sd25,
8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd14,
8'sd0,
-8'sd1,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd46,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd64,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22
},
{8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd46,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd62,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd69,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd93,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
-8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
-8'sd56,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd65,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd74,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
-8'sd70,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
-8'sd43,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd57,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd83,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd68,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd48,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd59,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd57,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
-8'sd60,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
-8'sd58,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
-8'sd26,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
-8'sd28,
8'sd24,
8'sd17,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd50,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
-8'sd15,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd39,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd58,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd80,
-8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd58,
-8'sd71,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
-8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd56,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd5,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
-8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd64,
-8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
-8'sd6,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
-8'sd20,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd79,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd83,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
-8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44
},
{8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd128,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
-8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd26,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd65,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd64,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd3,
8'sd0,
8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd56,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd37,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd99,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
-8'sd45,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
-8'sd4,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd33,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd90,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
-8'sd46,
-8'sd3,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd58,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd56,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd58,
8'sd0,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0
},
{8'sd0,
-8'sd61,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
-8'sd35,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
-8'sd22,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd58,
8'sd0,
-8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
-8'sd23,
8'sd71,
8'sd0,
-8'sd24,
8'sd0,
8'sd11,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
-8'sd80,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
-8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
-8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd46,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd57,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
-8'sd31,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd81,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd61,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd37,
-8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd36,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
-8'sd68,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd61,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd37,
8'sd95,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd0,
8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
-8'sd54,
8'sd0,
8'sd0,
-8'sd69,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
-8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd46,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd74,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
-8'sd22,
8'sd0,
8'sd0,
-8'sd18,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd63,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd56,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd52,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd76,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd7,
8'sd0,
8'sd57,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd56,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd87,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd57,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd57,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd69,
8'sd38,
8'sd4,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd59,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd58,
8'sd0,
8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd23,
8'sd0,
8'sd2,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd6,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
-8'sd51,
8'sd0,
8'sd0,
8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
-8'sd54,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd53,
-8'sd24,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd63,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd56,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
-8'sd58,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd12,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd71,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd62,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd59,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd7,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd39,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd60,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd13,
8'sd0,
8'sd19,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd82,
8'sd0,
8'sd0,
-8'sd20,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
-8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
8'sd25,
8'sd0,
8'sd25,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd44,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
-8'sd22,
-8'sd19,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd44,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0
},
{-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
-8'sd41,
-8'sd14,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd62,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd66,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
-8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd14,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd5,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd72,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd66,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd25,
8'sd18,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd59,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd69,
8'sd0,
8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd56,
8'sd0,
8'sd101,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd59,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd33,
8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd23,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd53,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
-8'sd31,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
-8'sd77,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd51,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd84,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd11,
8'sd50,
8'sd0,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
-8'sd42,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd53,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
-8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
-8'sd56,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
-8'sd7,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd64,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
-8'sd27,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd63,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
-8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd55,
8'sd13,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
-8'sd8,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd46,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd56,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd48,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
-8'sd10,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd49,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd59,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd60,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd56,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd35,
-8'sd9,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
-8'sd29,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd78,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd14,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd49
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
-8'sd26,
8'sd0,
-8'sd7,
8'sd0,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd56,
8'sd0,
8'sd5,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd33,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
-8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd65,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
-8'sd8,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd58,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd58,
8'sd0,
8'sd73,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd94,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
-8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd66,
8'sd0,
-8'sd20,
8'sd0,
-8'sd44,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
-8'sd76,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd52,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd7,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
-8'sd63,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd55,
-8'sd33,
8'sd0,
8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd59,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd58,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
-8'sd68,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
-8'sd8,
8'sd0,
8'sd59,
8'sd0,
8'sd0,
8'sd44,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd59
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
-8'sd4,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd82,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd48,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd70,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd62,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
-8'sd21,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd65,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd45,
8'sd0,
8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd45,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
-8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd65,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd29,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd69,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd55,
8'sd0,
-8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd46,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd59,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
-8'sd79,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd55,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd57,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd18,
8'sd0
},
{8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd52,
8'sd0,
8'sd0,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd20,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd64,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
-8'sd18,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd74,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd59,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd57,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd76,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
-8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd56,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
-8'sd29,
8'sd0,
8'sd0,
8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd50,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd58,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd80,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd49,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
-8'sd4
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd52,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
-8'sd64,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd83,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd37,
8'sd0,
-8'sd3,
8'sd0,
8'sd55,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd12,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd16,
-8'sd51,
8'sd28,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd67,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
-8'sd48,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd62,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd31,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd7,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd50,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
-8'sd55,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd53,
8'sd64,
8'sd0,
8'sd32,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
-8'sd69,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd58,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd30,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd65,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd33,
8'sd0,
8'sd7,
8'sd0,
-8'sd92,
8'sd0,
8'sd33,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd95,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
-8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd75,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd69,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd48,
8'sd0,
8'sd0,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd88,
8'sd0,
8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd2,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd66,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd47,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd89,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd56,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
-8'sd69,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
-8'sd58,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
-8'sd42,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
-8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
-8'sd19,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
-8'sd60,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd82,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd33,
8'sd0,
8'sd65,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd51,
-8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd30,
8'sd0,
8'sd58,
8'sd0,
8'sd0,
8'sd0,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd62,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{-8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd22
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd56,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
-8'sd33,
8'sd0,
8'sd0,
8'sd0,
-8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
-8'sd4,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd15,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd60,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd8,
-8'sd62,
8'sd0,
8'sd0,
8'sd0,
8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd46,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
-8'sd11,
8'sd0,
-8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
-8'sd10,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd62,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd44,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd8,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
-8'sd75,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd65,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd61,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd77,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd21,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd36,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd49,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd47,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
-8'sd5,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd55,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd48,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
-8'sd57,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
-8'sd6,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd81,
8'sd59,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd77,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd62,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd72,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd7,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd37,
8'sd0,
8'sd0,
-8'sd30,
8'sd28,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd28,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd38,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0
},
{8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd48,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd47,
8'sd12,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd18,
8'sd0,
8'sd58,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd3,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
-8'sd18,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd30,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd0,
8'sd0,
8'sd29,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{-8'sd2,
8'sd0,
8'sd0,
8'sd5,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd50,
8'sd0,
8'sd0,
8'sd53,
8'sd0,
-8'sd32,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
-8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd42,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
-8'sd80,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd53,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd1,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd0,
-8'sd39,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd45,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
-8'sd2,
8'sd0,
8'sd17,
-8'sd61,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd23,
8'sd0,
8'sd0,
8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd43,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd52,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd58,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd56,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd14,
-8'sd16,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd23,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd50,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd60,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd17,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd32,
8'sd7,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd63,
-8'sd1,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd55,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd16,
-8'sd51,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd36,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd65,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd9,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd13,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd41,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd15,
8'sd0,
8'sd17,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd12,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd33,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
-8'sd22,
8'sd0,
8'sd0
},
{8'sd72,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd64,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd25,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd40,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd16,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd35,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd83,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd37,
8'sd0,
8'sd0,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd60,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd54,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd36,
8'sd0,
8'sd0,
8'sd26,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd36,
8'sd0,
8'sd0,
8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd15,
8'sd0,
8'sd0,
8'sd0,
8'sd59,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd31,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd8,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd34,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd77,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd61,
8'sd0,
8'sd0,
8'sd0,
8'sd10,
8'sd0,
-8'sd32,
8'sd0,
8'sd65,
8'sd0,
-8'sd27,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd66,
8'sd18,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd20,
8'sd0,
8'sd10,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd4,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd5,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd90,
8'sd0,
8'sd0,
8'sd39,
8'sd0,
8'sd0,
-8'sd14,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd40,
8'sd0,
8'sd0,
8'sd0
},
{8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd19,
-8'sd57,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd1,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd9,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd24,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd2,
8'sd0,
8'sd0,
8'sd0,
8'sd22,
8'sd6,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd19,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd36,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd28,
8'sd0,
8'sd0,
8'sd0,
-8'sd26,
8'sd0,
8'sd0,
8'sd0,
-8'sd22,
8'sd46,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd11,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd2,
8'sd0,
8'sd0,
-8'sd20,
8'sd0,
-8'sd30,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
-8'sd21,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0,
8'sd0
}
};
// Output layer
reg signed [7:0] output_weight [0: num_reservoir_neurons-1];initial {
	output_weight[0],
output_weight[1],
output_weight[2],
output_weight[3],
output_weight[4],
output_weight[5],
output_weight[6],
output_weight[7],
output_weight[8],
output_weight[9],
output_weight[10],
output_weight[11],
output_weight[12],
output_weight[13],
output_weight[14],
output_weight[15],
output_weight[16],
output_weight[17],
output_weight[18],
output_weight[19],
output_weight[20],
output_weight[21],
output_weight[22],
output_weight[23],
output_weight[24],
output_weight[25],
output_weight[26],
output_weight[27],
output_weight[28],
output_weight[29],
output_weight[30],
output_weight[31],
output_weight[32],
output_weight[33],
output_weight[34],
output_weight[35],
output_weight[36],
output_weight[37],
output_weight[38],
output_weight[39],
output_weight[40],
output_weight[41],
output_weight[42],
output_weight[43],
output_weight[44],
output_weight[45],
output_weight[46],
output_weight[47],
output_weight[48],
output_weight[49],
output_weight[50],
output_weight[51],
output_weight[52],
output_weight[53],
output_weight[54],
output_weight[55],
output_weight[56],
output_weight[57],
output_weight[58],
output_weight[59],
output_weight[60],
output_weight[61],
output_weight[62],
output_weight[63],
output_weight[64],
output_weight[65],
output_weight[66],
output_weight[67],
output_weight[68],
output_weight[69],
output_weight[70],
output_weight[71],
output_weight[72],
output_weight[73],
output_weight[74],
output_weight[75],
output_weight[76],
output_weight[77],
output_weight[78],
output_weight[79],
output_weight[80],
output_weight[81],
output_weight[82],
output_weight[83],
output_weight[84],
output_weight[85],
output_weight[86],
output_weight[87],
output_weight[88],
output_weight[89],
output_weight[90],
output_weight[91],
output_weight[92],
output_weight[93],
output_weight[94],
output_weight[95],
output_weight[96],
output_weight[97],
output_weight[98],
output_weight[99],
output_weight[100],
output_weight[101],
output_weight[102],
output_weight[103],
output_weight[104],
output_weight[105],
output_weight[106],
output_weight[107],
output_weight[108],
output_weight[109],
output_weight[110],
output_weight[111],
output_weight[112],
output_weight[113],
output_weight[114],
output_weight[115],
output_weight[116],
output_weight[117],
output_weight[118],
output_weight[119],
output_weight[120],
output_weight[121],
output_weight[122],
output_weight[123],
output_weight[124],
output_weight[125],
output_weight[126],
output_weight[127],
output_weight[128],
output_weight[129],
output_weight[130],
output_weight[131],
output_weight[132],
output_weight[133],
output_weight[134],
output_weight[135],
output_weight[136],
output_weight[137],
output_weight[138],
output_weight[139],
output_weight[140],
output_weight[141],
output_weight[142],
output_weight[143],
output_weight[144],
output_weight[145],
output_weight[146],
output_weight[147],
output_weight[148],
output_weight[149],
output_weight[150],
output_weight[151],
output_weight[152],
output_weight[153],
output_weight[154],
output_weight[155],
output_weight[156],
output_weight[157],
output_weight[158],
output_weight[159],
output_weight[160],
output_weight[161],
output_weight[162],
output_weight[163],
output_weight[164],
output_weight[165],
output_weight[166],
output_weight[167],
output_weight[168],
output_weight[169],
output_weight[170],
output_weight[171],
output_weight[172],
output_weight[173],
output_weight[174],
output_weight[175],
output_weight[176],
output_weight[177],
output_weight[178],
output_weight[179],
output_weight[180],
output_weight[181],
output_weight[182],
output_weight[183],
output_weight[184],
output_weight[185],
output_weight[186],
output_weight[187],
output_weight[188],
output_weight[189],
output_weight[190],
output_weight[191],
output_weight[192],
output_weight[193],
output_weight[194],
output_weight[195],
output_weight[196],
output_weight[197],
output_weight[198],
output_weight[199]
} = {
-8'sd3,
8'sd5,
8'sd4,
8'sd2,
8'sd0,
-8'sd2,
8'sd2,
-8'sd6,
8'sd0,
8'sd4,
8'sd2,
8'sd5,
8'sd2,
-8'sd3,
8'sd3,
8'sd17,
-8'sd11,
-8'sd2,
8'sd3,
8'sd15,
8'sd4,
-8'sd1,
8'sd3,
8'sd8,
8'sd2,
8'sd50,
8'sd6,
8'sd6,
8'sd5,
8'sd0,
-8'sd2,
8'sd8,
-8'sd5,
8'sd2,
8'sd4,
8'sd7,
-8'sd2,
8'sd3,
-8'sd6,
-8'sd6,
8'sd2,
8'sd0,
8'sd9,
-8'sd1,
8'sd2,
-8'sd4,
-8'sd7,
8'sd3,
-8'sd2,
8'sd0,
8'sd6,
8'sd9,
-8'sd3,
8'sd7,
8'sd0,
-8'sd5,
8'sd2,
8'sd7,
-8'sd3,
8'sd3,
8'sd0,
8'sd1,
-8'sd2,
8'sd8,
-8'sd2,
8'sd5,
8'sd2,
8'sd1,
8'sd0,
8'sd1,
-8'sd6,
8'sd2,
-8'sd5,
-8'sd5,
8'sd5,
8'sd1,
-8'sd2,
-8'sd4,
-8'sd1,
-8'sd2,
8'sd7,
8'sd1,
-8'sd1,
-8'sd4,
-8'sd8,
8'sd1,
8'sd4,
-8'sd8,
8'sd1,
8'sd12,
8'sd8,
-8'sd5,
8'sd5,
-8'sd1,
8'sd0,
-8'sd1,
8'sd5,
-8'sd1,
8'sd4,
8'sd0,
-8'sd5,
8'sd2,
-8'sd2,
-8'sd2,
8'sd0,
8'sd5,
8'sd3,
8'sd1,
8'sd9,
-8'sd4,
8'sd0,
8'sd3,
-8'sd6,
-8'sd6,
-8'sd3,
-8'sd6,
8'sd1,
8'sd5,
8'sd6,
-8'sd1,
-8'sd5,
-8'sd3,
8'sd5,
8'sd3,
-8'sd2,
-8'sd1,
8'sd6,
8'sd2,
8'sd3,
-8'sd2,
8'sd0,
8'sd1,
8'sd1,
8'sd3,
8'sd6,
-8'sd1,
8'sd0,
8'sd5,
-8'sd4,
-8'sd1,
-8'sd1,
8'sd4,
-8'sd2,
-8'sd1,
-8'sd4,
-8'sd1,
-8'sd5,
8'sd7,
8'sd2,
8'sd10,
-8'sd3,
-8'sd2,
-8'sd2,
-8'sd3,
-8'sd2,
-8'sd127,
-8'sd8,
-8'sd2,
-8'sd4,
8'sd5,
-8'sd4,
-8'sd1,
-8'sd2,
8'sd0,
-8'sd7,
8'sd5,
-8'sd5,
-8'sd2,
8'sd0,
8'sd2,
8'sd5,
8'sd4,
8'sd2,
8'sd6,
-8'sd8,
8'sd3,
8'sd3,
8'sd6,
-8'sd11,
-8'sd8,
8'sd3,
-8'sd8,
8'sd9,
-8'sd3,
8'sd3,
8'sd7,
-8'sd4,
8'sd2,
-8'sd3,
8'sd2,
-8'sd2,
8'sd2,
8'sd1,
-8'sd3,
-8'sd1,
-8'sd1,
-8'sd2,
-8'sd2,
-8'sd5,
-8'sd5
};"
  // Scaling factors and zero point
  reg signed [31:0] scale = 32'b00000000000000010101101110001010;

  reg signed [31:0] input_sum_parallel [0: num_reservoir_neurons-1];
  reg signed [31:0] reservoir_sum_parallel [0: num_reservoir_neurons-1];
  reg signed [31:0] output_sum;
  integer i,j,k,x,y,t,m,n,p,q;

  reg signed [31:0] reg_input [0: num_reservoir_neurons-1];
  reg signed [31:0] reg_reservoir [0: num_reservoir_neurons-1];
  // ESN logic
  always @(posedge clk) begin

      for (i = 0; i < num_reservoir_neurons; i = i + 1) begin
        input_sum_parallel[i] = input_data * input_weight[i];
        reservoir_sum_parallel[i]= 0;
      end

      for (j = 0; j < num_reservoir_neurons; j = j + 1) begin
        for (k = 0; k < num_reservoir_neurons; k = k + 1) begin
          reservoir_sum_parallel[j] = reservoir_sum_parallel[j] + (reservoir_state[k] * reservoir_weight[k][j]);
        end
      end


      for (m = 0; m < num_reservoir_neurons; m = m + 1) begin
          reg_input[m] = 0;
          if (input_sum_parallel[m] < a_scaled) begin
              reg_input[m] = a_scaled;
          end
          else if (input_sum_parallel[m] > b_scaled) begin
              reg_input[m] = b_scaled;
          end
          else begin
              reg_input[m] = input_sum_parallel[m];
          end
      end

      for (p = 0; p < num_reservoir_neurons; p = p + 1) begin
          reg_reservoir[p] = 0;
          if (reservoir_sum_parallel[p] < c_scaled) begin
              reg_reservoir[p] = c_scaled;
          end
          else if (reservoir_sum_parallel[p] > d_scaled) begin
              reg_reservoir[p] = d_scaled;
          end
          else begin
              reg_reservoir[p] = reservoir_sum_parallel[p];
          end
      end

      for (k = 0; k < num_reservoir_neurons; k = k + 1) begin
          reg_input[j]=reg_input[j]+16'd1628;
          reg_input[k] <= reg_input[k] >> 8;
          reg_reservoir[k]=reg_reservoir[k]+16'd17641;
          reg_reservoir[k]<= reg_reservoir[k] >> 8;
      end

      for (y = 0; y < num_reservoir_neurons; y = y + 1) begin
          reservoir_state[y] <= reg_reservoir[y] + reg_input[y];

      end

      // Output calculation
       // Wider format for accumulation
      output_sum = 0;



      for (t = 0; t < num_reservoir_neurons; t = t + 1) begin
        output_sum = output_sum +(reservoir_state[t] * output_weight[t]);
      end




    end
    //assign output_data = output_sum * scale;
    assign output_data = output_sum ;
endmodule
